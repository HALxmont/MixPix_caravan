magic
tech sky130B
magscale 1 2
timestamp 1667049779
<< metal1 >>
rect 49694 702992 49700 703044
rect 49752 703032 49758 703044
rect 50890 703032 50896 703044
rect 49752 703004 50896 703032
rect 49752 702992 49758 703004
rect 50890 702992 50896 703004
rect 50948 702992 50954 703044
rect 69014 702992 69020 703044
rect 69072 703032 69078 703044
rect 70210 703032 70216 703044
rect 69072 703004 70216 703032
rect 69072 702992 69078 703004
rect 70210 702992 70216 703004
rect 70268 702992 70274 703044
rect 309134 702992 309140 703044
rect 309192 703032 309198 703044
rect 310422 703032 310428 703044
rect 309192 703004 310428 703032
rect 309192 702992 309198 703004
rect 310422 702992 310428 703004
rect 310480 702992 310486 703044
rect 328454 702992 328460 703044
rect 328512 703032 328518 703044
rect 329742 703032 329748 703044
rect 328512 703004 329748 703032
rect 328512 702992 328518 703004
rect 329742 702992 329748 703004
rect 329800 702992 329806 703044
rect 347774 702992 347780 703044
rect 347832 703032 347838 703044
rect 349062 703032 349068 703044
rect 347832 703004 349068 703032
rect 347832 702992 347838 703004
rect 349062 702992 349068 703004
rect 349120 702992 349126 703044
rect 358814 702992 358820 703044
rect 358872 703032 358878 703044
rect 360010 703032 360016 703044
rect 358872 703004 360016 703032
rect 358872 702992 358878 703004
rect 360010 702992 360016 703004
rect 360068 702992 360074 703044
rect 378134 702992 378140 703044
rect 378192 703032 378198 703044
rect 379330 703032 379336 703044
rect 378192 703004 379336 703032
rect 378192 702992 378198 703004
rect 379330 702992 379336 703004
rect 379388 702992 379394 703044
rect 576118 702448 576124 702500
rect 576176 702488 576182 702500
rect 580166 702488 580172 702500
rect 576176 702460 580172 702488
rect 576176 702448 576182 702460
rect 580166 702448 580172 702460
rect 580224 702448 580230 702500
rect 3050 701020 3056 701072
rect 3108 701060 3114 701072
rect 98638 701060 98644 701072
rect 3108 701032 98644 701060
rect 3108 701020 3114 701032
rect 98638 701020 98644 701032
rect 98696 701020 98702 701072
rect 184842 700612 184848 700664
rect 184900 700652 184906 700664
rect 195974 700652 195980 700664
rect 184900 700624 195980 700652
rect 184900 700612 184906 700624
rect 195974 700612 195980 700624
rect 196032 700612 196038 700664
rect 188062 700544 188068 700596
rect 188120 700584 188126 700596
rect 200114 700584 200120 700596
rect 188120 700556 200120 700584
rect 188120 700544 188126 700556
rect 200114 700544 200120 700556
rect 200172 700544 200178 700596
rect 66346 700476 66352 700528
rect 66404 700516 66410 700528
rect 78030 700516 78036 700528
rect 66404 700488 78036 700516
rect 66404 700476 66410 700488
rect 78030 700476 78036 700488
rect 78088 700476 78094 700528
rect 115842 700476 115848 700528
rect 115900 700516 115906 700528
rect 123662 700516 123668 700528
rect 115900 700488 123668 700516
rect 115900 700476 115906 700488
rect 123662 700476 123668 700488
rect 123720 700476 123726 700528
rect 177114 700476 177120 700528
rect 177172 700516 177178 700528
rect 194686 700516 194692 700528
rect 177172 700488 194692 700516
rect 177172 700476 177178 700488
rect 194686 700476 194692 700488
rect 194744 700476 194750 700528
rect 19978 700408 19984 700460
rect 20036 700448 20042 700460
rect 31018 700448 31024 700460
rect 20036 700420 31024 700448
rect 20036 700408 20042 700420
rect 31018 700408 31024 700420
rect 31076 700408 31082 700460
rect 77294 700408 77300 700460
rect 77352 700448 77358 700460
rect 116026 700448 116032 700460
rect 77352 700420 116032 700448
rect 77352 700408 77358 700420
rect 116026 700408 116032 700420
rect 116084 700408 116090 700460
rect 169386 700408 169392 700460
rect 169444 700448 169450 700460
rect 191834 700448 191840 700460
rect 169444 700420 191840 700448
rect 169444 700408 169450 700420
rect 191834 700408 191840 700420
rect 191892 700408 191898 700460
rect 194502 700408 194508 700460
rect 194560 700448 194566 700460
rect 287882 700448 287888 700460
rect 194560 700420 287888 700448
rect 194560 700408 194566 700420
rect 287882 700408 287888 700420
rect 287940 700408 287946 700460
rect 16114 700340 16120 700392
rect 16172 700380 16178 700392
rect 77938 700380 77944 700392
rect 16172 700352 77944 700380
rect 16172 700340 16178 700352
rect 77938 700340 77944 700352
rect 77996 700340 78002 700392
rect 117222 700340 117228 700392
rect 117280 700380 117286 700392
rect 127526 700380 127532 700392
rect 117280 700352 127532 700380
rect 117280 700340 117286 700352
rect 127526 700340 127532 700352
rect 127584 700340 127590 700392
rect 165522 700340 165528 700392
rect 165580 700380 165586 700392
rect 193214 700380 193220 700392
rect 165580 700352 193220 700380
rect 165580 700340 165586 700352
rect 193214 700340 193220 700352
rect 193272 700340 193278 700392
rect 199378 700340 199384 700392
rect 199436 700380 199442 700392
rect 394786 700380 394792 700392
rect 199436 700352 394792 700380
rect 199436 700340 199442 700352
rect 394786 700340 394792 700352
rect 394844 700340 394850 700392
rect 548610 700340 548616 700392
rect 548668 700380 548674 700392
rect 570598 700380 570604 700392
rect 548668 700352 570604 700380
rect 548668 700340 548674 700352
rect 570598 700340 570604 700352
rect 570656 700340 570662 700392
rect 31570 700272 31576 700324
rect 31628 700312 31634 700324
rect 113174 700312 113180 700324
rect 31628 700284 113180 700312
rect 31628 700272 31634 700284
rect 113174 700272 113180 700284
rect 113232 700272 113238 700324
rect 121270 700272 121276 700324
rect 121328 700312 121334 700324
rect 157794 700312 157800 700324
rect 121328 700284 157800 700312
rect 121328 700272 121334 700284
rect 157794 700272 157800 700284
rect 157852 700272 157858 700324
rect 189718 700272 189724 700324
rect 189776 700312 189782 700324
rect 551278 700312 551284 700324
rect 189776 700284 551284 700312
rect 189776 700272 189782 700284
rect 551278 700272 551284 700284
rect 551336 700272 551342 700324
rect 556798 700272 556804 700324
rect 556856 700312 556862 700324
rect 574462 700312 574468 700324
rect 556856 700284 574468 700312
rect 556856 700272 556862 700284
rect 574462 700272 574468 700284
rect 574520 700272 574526 700324
rect 180978 700068 180984 700120
rect 181036 700108 181042 700120
rect 189442 700108 189448 700120
rect 181036 700080 189448 700108
rect 181036 700068 181042 700080
rect 189442 700068 189448 700080
rect 189500 700068 189506 700120
rect 115934 699796 115940 699848
rect 115992 699836 115998 699848
rect 117958 699836 117964 699848
rect 115992 699808 117964 699836
rect 115992 699796 115998 699808
rect 117958 699796 117964 699808
rect 118016 699796 118022 699848
rect 119798 699660 119804 699712
rect 119856 699700 119862 699712
rect 120718 699700 120724 699712
rect 119856 699672 120724 699700
rect 119856 699660 119862 699672
rect 120718 699660 120724 699672
rect 120776 699660 120782 699712
rect 199654 699660 199660 699712
rect 199712 699700 199718 699712
rect 201494 699700 201500 699712
rect 199712 699672 201500 699700
rect 199712 699660 199718 699672
rect 201494 699660 201500 699672
rect 201552 699660 201558 699712
rect 220078 699660 220084 699712
rect 220136 699700 220142 699712
rect 222838 699700 222844 699712
rect 220136 699672 222844 699700
rect 220136 699660 220142 699672
rect 222838 699660 222844 699672
rect 222896 699660 222902 699712
rect 224218 699660 224224 699712
rect 224276 699700 224282 699712
rect 226702 699700 226708 699712
rect 224276 699672 226708 699700
rect 224276 699660 224282 699672
rect 226702 699660 226708 699672
rect 226760 699660 226766 699712
rect 242158 699660 242164 699712
rect 242216 699700 242222 699712
rect 245378 699700 245384 699712
rect 242216 699672 245384 699700
rect 242216 699660 242222 699672
rect 245378 699660 245384 699672
rect 245436 699660 245442 699712
rect 269758 699660 269764 699712
rect 269816 699700 269822 699712
rect 272426 699700 272432 699712
rect 269816 699672 272432 699700
rect 269816 699660 269822 699672
rect 272426 699660 272432 699672
rect 272484 699660 272490 699712
rect 278038 699660 278044 699712
rect 278096 699700 278102 699712
rect 280154 699700 280160 699712
rect 278096 699672 280160 699700
rect 278096 699660 278102 699672
rect 280154 699660 280160 699672
rect 280212 699660 280218 699712
rect 323578 699660 323584 699712
rect 323636 699700 323642 699712
rect 325878 699700 325884 699712
rect 323636 699672 325884 699700
rect 323636 699660 323642 699672
rect 325878 699660 325884 699672
rect 325936 699660 325942 699712
rect 374638 699660 374644 699712
rect 374696 699700 374702 699712
rect 375466 699700 375472 699712
rect 374696 699672 375472 699700
rect 374696 699660 374702 699672
rect 375466 699660 375472 699672
rect 375524 699660 375530 699712
rect 395338 699660 395344 699712
rect 395396 699700 395402 699712
rect 398650 699700 398656 699712
rect 395396 699672 398656 699700
rect 395396 699660 395402 699672
rect 398650 699660 398656 699672
rect 398708 699660 398714 699712
rect 400858 699660 400864 699712
rect 400916 699700 400922 699712
rect 402514 699700 402520 699712
rect 400916 699672 402520 699700
rect 400916 699660 400922 699672
rect 402514 699660 402520 699672
rect 402572 699660 402578 699712
rect 445018 699660 445024 699712
rect 445076 699700 445082 699712
rect 448238 699700 448244 699712
rect 445076 699672 448244 699700
rect 445076 699660 445082 699672
rect 448238 699660 448244 699672
rect 448296 699660 448302 699712
rect 449158 699660 449164 699712
rect 449216 699700 449222 699712
rect 452102 699700 452108 699712
rect 449216 699672 452108 699700
rect 449216 699660 449222 699672
rect 452102 699660 452108 699672
rect 452160 699660 452166 699712
rect 472618 699660 472624 699712
rect 472676 699700 472682 699712
rect 474642 699700 474648 699712
rect 472676 699672 474648 699700
rect 472676 699660 472682 699672
rect 474642 699660 474648 699672
rect 474700 699660 474706 699712
rect 494698 699660 494704 699712
rect 494756 699700 494762 699712
rect 497826 699700 497832 699712
rect 494756 699672 497832 699700
rect 494756 699660 494762 699672
rect 497826 699660 497832 699672
rect 497884 699660 497890 699712
rect 498838 699660 498844 699712
rect 498896 699700 498902 699712
rect 501690 699700 501696 699712
rect 498896 699672 501696 699700
rect 498896 699660 498902 699672
rect 501690 699660 501696 699672
rect 501748 699660 501754 699712
rect 502978 699660 502984 699712
rect 503036 699700 503042 699712
rect 505554 699700 505560 699712
rect 503036 699672 505560 699700
rect 503036 699660 503042 699672
rect 505554 699660 505560 699672
rect 505612 699660 505618 699712
rect 552658 699660 552664 699712
rect 552716 699700 552722 699712
rect 555142 699700 555148 699712
rect 552716 699672 555148 699700
rect 552716 699660 552722 699672
rect 555142 699660 555148 699672
rect 555200 699660 555206 699712
rect 570598 698300 570604 698352
rect 570656 698340 570662 698352
rect 580166 698340 580172 698352
rect 570656 698312 580172 698340
rect 570656 698300 570662 698312
rect 580166 698300 580172 698312
rect 580224 698300 580230 698352
rect 144914 697552 144920 697604
rect 144972 697592 144978 697604
rect 146202 697592 146208 697604
rect 144972 697564 146208 697592
rect 144972 697552 144978 697564
rect 146202 697552 146208 697564
rect 146260 697552 146266 697604
rect 492674 697552 492680 697604
rect 492732 697592 492738 697604
rect 493962 697592 493968 697604
rect 492732 697564 493968 697592
rect 492732 697552 492738 697564
rect 493962 697552 493968 697564
rect 494020 697552 494026 697604
rect 511994 697552 512000 697604
rect 512052 697592 512058 697604
rect 513282 697592 513288 697604
rect 512052 697564 513288 697592
rect 512052 697552 512058 697564
rect 513282 697552 513288 697564
rect 513340 697552 513346 697604
rect 544378 694152 544384 694204
rect 544436 694192 544442 694204
rect 580166 694192 580172 694204
rect 544436 694164 580172 694192
rect 544436 694152 544442 694164
rect 580166 694152 580172 694164
rect 580224 694152 580230 694204
rect 3142 692792 3148 692844
rect 3200 692832 3206 692844
rect 88978 692832 88984 692844
rect 3200 692804 88984 692832
rect 3200 692792 3206 692804
rect 88978 692792 88984 692804
rect 89036 692792 89042 692844
rect 3418 688644 3424 688696
rect 3476 688684 3482 688696
rect 89070 688684 89076 688696
rect 3476 688656 89076 688684
rect 3476 688644 3482 688656
rect 89070 688644 89076 688656
rect 89128 688644 89134 688696
rect 548518 685856 548524 685908
rect 548576 685896 548582 685908
rect 579798 685896 579804 685908
rect 548576 685868 579804 685896
rect 548576 685856 548582 685868
rect 579798 685856 579804 685868
rect 579856 685856 579862 685908
rect 3142 684496 3148 684548
rect 3200 684536 3206 684548
rect 181438 684536 181444 684548
rect 3200 684508 181444 684536
rect 3200 684496 3206 684508
rect 181438 684496 181444 684508
rect 181496 684496 181502 684548
rect 3418 680348 3424 680400
rect 3476 680388 3482 680400
rect 94498 680388 94504 680400
rect 3476 680360 94504 680388
rect 3476 680348 3482 680360
rect 94498 680348 94504 680360
rect 94556 680348 94562 680400
rect 576210 677560 576216 677612
rect 576268 677600 576274 677612
rect 580166 677600 580172 677612
rect 576268 677572 580172 677600
rect 576268 677560 576274 677572
rect 580166 677560 580172 677572
rect 580224 677560 580230 677612
rect 3234 672052 3240 672104
rect 3292 672092 3298 672104
rect 105538 672092 105544 672104
rect 3292 672064 105544 672092
rect 3292 672052 3298 672064
rect 105538 672052 105544 672064
rect 105596 672052 105602 672104
rect 556890 669332 556896 669384
rect 556948 669372 556954 669384
rect 580166 669372 580172 669384
rect 556948 669344 580172 669372
rect 556948 669332 556954 669344
rect 580166 669332 580172 669344
rect 580224 669332 580230 669384
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 84838 667944 84844 667956
rect 3476 667916 84844 667944
rect 3476 667904 3482 667916
rect 84838 667904 84844 667916
rect 84896 667904 84902 667956
rect 202138 665184 202144 665236
rect 202196 665224 202202 665236
rect 580166 665224 580172 665236
rect 202196 665196 580172 665224
rect 202196 665184 202202 665196
rect 580166 665184 580172 665196
rect 580224 665184 580230 665236
rect 3234 663756 3240 663808
rect 3292 663796 3298 663808
rect 111886 663796 111892 663808
rect 3292 663768 111892 663796
rect 3292 663756 3298 663768
rect 111886 663756 111892 663768
rect 111944 663756 111950 663808
rect 3418 661036 3424 661088
rect 3476 661076 3482 661088
rect 80698 661076 80704 661088
rect 3476 661048 80704 661076
rect 3476 661036 3482 661048
rect 80698 661036 80704 661048
rect 80756 661036 80762 661088
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 111058 652780 111064 652792
rect 3108 652752 111064 652780
rect 3108 652740 3114 652752
rect 111058 652740 111064 652752
rect 111116 652740 111122 652792
rect 196618 648592 196624 648644
rect 196676 648632 196682 648644
rect 579982 648632 579988 648644
rect 196676 648604 579988 648632
rect 196676 648592 196682 648604
rect 579982 648592 579988 648604
rect 580040 648592 580046 648644
rect 3418 644444 3424 644496
rect 3476 644484 3482 644496
rect 98730 644484 98736 644496
rect 3476 644456 98736 644484
rect 3476 644444 3482 644456
rect 98730 644444 98736 644456
rect 98788 644444 98794 644496
rect 566458 644444 566464 644496
rect 566516 644484 566522 644496
rect 580166 644484 580172 644496
rect 566516 644456 580172 644484
rect 566516 644444 566522 644456
rect 580166 644444 580172 644456
rect 580224 644444 580230 644496
rect 567838 633428 567844 633480
rect 567896 633468 567902 633480
rect 580166 633468 580172 633480
rect 567896 633440 580172 633468
rect 567896 633428 567902 633440
rect 580166 633428 580172 633440
rect 580224 633428 580230 633480
rect 552750 629280 552756 629332
rect 552808 629320 552814 629332
rect 580166 629320 580172 629332
rect 552808 629292 580172 629320
rect 552808 629280 552814 629292
rect 580166 629280 580172 629292
rect 580224 629280 580230 629332
rect 3418 627920 3424 627972
rect 3476 627960 3482 627972
rect 95878 627960 95884 627972
rect 3476 627932 95884 627960
rect 3476 627920 3482 627932
rect 95878 627920 95884 627932
rect 95936 627920 95942 627972
rect 577498 625404 577504 625456
rect 577556 625444 577562 625456
rect 580534 625444 580540 625456
rect 577556 625416 580540 625444
rect 577556 625404 577562 625416
rect 580534 625404 580540 625416
rect 580592 625404 580598 625456
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 128354 623812 128360 623824
rect 3292 623784 128360 623812
rect 3292 623772 3298 623784
rect 128354 623772 128360 623784
rect 128412 623772 128418 623824
rect 3418 619624 3424 619676
rect 3476 619664 3482 619676
rect 106918 619664 106924 619676
rect 3476 619636 106924 619664
rect 3476 619624 3482 619636
rect 106918 619624 106924 619636
rect 106976 619624 106982 619676
rect 3234 615476 3240 615528
rect 3292 615516 3298 615528
rect 98822 615516 98828 615528
rect 3292 615488 98828 615516
rect 3292 615476 3298 615488
rect 98822 615476 98828 615488
rect 98880 615476 98886 615528
rect 3418 612756 3424 612808
rect 3476 612796 3482 612808
rect 97258 612796 97264 612808
rect 3476 612768 97264 612796
rect 3476 612756 3482 612768
rect 97258 612756 97264 612768
rect 97316 612756 97322 612808
rect 3418 608608 3424 608660
rect 3476 608648 3482 608660
rect 125686 608648 125692 608660
rect 3476 608620 125692 608648
rect 3476 608608 3482 608620
rect 125686 608608 125692 608620
rect 125744 608608 125750 608660
rect 565078 608608 565084 608660
rect 565136 608648 565142 608660
rect 580166 608648 580172 608660
rect 565136 608620 580172 608648
rect 565136 608608 565142 608620
rect 580166 608608 580172 608620
rect 580224 608608 580230 608660
rect 3418 604460 3424 604512
rect 3476 604500 3482 604512
rect 102778 604500 102784 604512
rect 3476 604472 102784 604500
rect 3476 604460 3482 604472
rect 102778 604460 102784 604472
rect 102836 604460 102842 604512
rect 3418 600312 3424 600364
rect 3476 600352 3482 600364
rect 86218 600352 86224 600364
rect 3476 600324 86224 600352
rect 3476 600312 3482 600324
rect 86218 600312 86224 600324
rect 86276 600312 86282 600364
rect 3418 596164 3424 596216
rect 3476 596204 3482 596216
rect 101398 596204 101404 596216
rect 3476 596176 101404 596204
rect 3476 596164 3482 596176
rect 101398 596164 101404 596176
rect 101456 596164 101462 596216
rect 567930 596164 567936 596216
rect 567988 596204 567994 596216
rect 580166 596204 580172 596216
rect 567988 596176 580172 596204
rect 567988 596164 567994 596176
rect 580166 596164 580172 596176
rect 580224 596164 580230 596216
rect 197998 592016 198004 592068
rect 198056 592056 198062 592068
rect 580166 592056 580172 592068
rect 198056 592028 580172 592056
rect 198056 592016 198062 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 3418 587868 3424 587920
rect 3476 587908 3482 587920
rect 95970 587908 95976 587920
rect 3476 587880 95976 587908
rect 3476 587868 3482 587880
rect 95970 587868 95976 587880
rect 96028 587868 96034 587920
rect 3418 583720 3424 583772
rect 3476 583760 3482 583772
rect 90358 583760 90364 583772
rect 3476 583732 90364 583760
rect 3476 583720 3482 583732
rect 90358 583720 90364 583732
rect 90416 583720 90422 583772
rect 574738 583720 574744 583772
rect 574796 583760 574802 583772
rect 580166 583760 580172 583772
rect 574796 583732 580172 583760
rect 574796 583720 574802 583732
rect 580166 583720 580172 583732
rect 580224 583720 580230 583772
rect 3418 579640 3424 579692
rect 3476 579680 3482 579692
rect 100018 579680 100024 579692
rect 3476 579652 100024 579680
rect 3476 579640 3482 579652
rect 100018 579640 100024 579652
rect 100076 579640 100082 579692
rect 3234 575492 3240 575544
rect 3292 575532 3298 575544
rect 102870 575532 102876 575544
rect 3292 575504 102876 575532
rect 3292 575492 3298 575504
rect 102870 575492 102876 575504
rect 102928 575492 102934 575544
rect 566642 572704 566648 572756
rect 566700 572744 566706 572756
rect 580166 572744 580172 572756
rect 566700 572716 580172 572744
rect 566700 572704 566706 572716
rect 580166 572704 580172 572716
rect 580224 572704 580230 572756
rect 3418 571344 3424 571396
rect 3476 571384 3482 571396
rect 90450 571384 90456 571396
rect 3476 571356 90456 571384
rect 3476 571344 3482 571356
rect 90450 571344 90456 571356
rect 90508 571344 90514 571396
rect 544470 568556 544476 568608
rect 544528 568596 544534 568608
rect 579706 568596 579712 568608
rect 544528 568568 579712 568596
rect 544528 568556 544534 568568
rect 579706 568556 579712 568568
rect 579764 568556 579770 568608
rect 3234 567196 3240 567248
rect 3292 567236 3298 567248
rect 91738 567236 91744 567248
rect 3292 567208 91744 567236
rect 3292 567196 3298 567208
rect 91738 567196 91744 567208
rect 91796 567196 91802 567248
rect 3418 564408 3424 564460
rect 3476 564448 3482 564460
rect 7558 564448 7564 564460
rect 3476 564420 7564 564448
rect 3476 564408 3482 564420
rect 7558 564408 7564 564420
rect 7616 564408 7622 564460
rect 571978 564408 571984 564460
rect 572036 564448 572042 564460
rect 580166 564448 580172 564460
rect 572036 564420 580172 564448
rect 572036 564408 572042 564420
rect 580166 564408 580172 564420
rect 580224 564408 580230 564460
rect 3418 560260 3424 560312
rect 3476 560300 3482 560312
rect 93118 560300 93124 560312
rect 3476 560272 93124 560300
rect 3476 560260 3482 560272
rect 93118 560260 93124 560272
rect 93176 560260 93182 560312
rect 200758 560260 200764 560312
rect 200816 560300 200822 560312
rect 579614 560300 579620 560312
rect 200816 560272 579620 560300
rect 200816 560260 200822 560272
rect 579614 560260 579620 560272
rect 579672 560260 579678 560312
rect 3418 556180 3424 556232
rect 3476 556220 3482 556232
rect 110414 556220 110420 556232
rect 3476 556192 110420 556220
rect 3476 556180 3482 556192
rect 110414 556180 110420 556192
rect 110472 556180 110478 556232
rect 3418 552032 3424 552084
rect 3476 552072 3482 552084
rect 112438 552072 112444 552084
rect 3476 552044 112444 552072
rect 3476 552032 3482 552044
rect 112438 552032 112444 552044
rect 112496 552032 112502 552084
rect 3234 547884 3240 547936
rect 3292 547924 3298 547936
rect 107010 547924 107016 547936
rect 3292 547896 107016 547924
rect 3292 547884 3298 547896
rect 107010 547884 107016 547896
rect 107068 547884 107074 547936
rect 193858 547884 193864 547936
rect 193916 547924 193922 547936
rect 580074 547924 580080 547936
rect 193916 547896 580080 547924
rect 193916 547884 193922 547896
rect 580074 547884 580080 547896
rect 580132 547884 580138 547936
rect 3326 543736 3332 543788
rect 3384 543776 3390 543788
rect 61378 543776 61384 543788
rect 3384 543748 61384 543776
rect 3384 543736 3390 543748
rect 61378 543736 61384 543748
rect 61436 543736 61442 543788
rect 554038 543736 554044 543788
rect 554096 543776 554102 543788
rect 580166 543776 580172 543788
rect 554096 543748 580172 543776
rect 554096 543736 554102 543748
rect 580166 543736 580172 543748
rect 580224 543736 580230 543788
rect 3418 539588 3424 539640
rect 3476 539628 3482 539640
rect 104158 539628 104164 539640
rect 3476 539600 104164 539628
rect 3476 539588 3482 539600
rect 104158 539588 104164 539600
rect 104216 539588 104222 539640
rect 570690 539588 570696 539640
rect 570748 539628 570754 539640
rect 579706 539628 579712 539640
rect 570748 539600 579712 539628
rect 570748 539588 570754 539600
rect 579706 539588 579712 539600
rect 579764 539588 579770 539640
rect 192478 535440 192484 535492
rect 192536 535480 192542 535492
rect 580166 535480 580172 535492
rect 192536 535452 580172 535480
rect 192536 535440 192542 535452
rect 580166 535440 580172 535452
rect 580224 535440 580230 535492
rect 3234 531292 3240 531344
rect 3292 531332 3298 531344
rect 94590 531332 94596 531344
rect 3292 531304 94596 531332
rect 3292 531292 3298 531304
rect 94590 531292 94596 531304
rect 94648 531292 94654 531344
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 10318 527184 10324 527196
rect 3476 527156 10324 527184
rect 3476 527144 3482 527156
rect 10318 527144 10324 527156
rect 10376 527144 10382 527196
rect 560938 527144 560944 527196
rect 560996 527184 561002 527196
rect 580166 527184 580172 527196
rect 560996 527156 580172 527184
rect 560996 527144 561002 527156
rect 580166 527144 580172 527156
rect 580224 527144 580230 527196
rect 3234 522996 3240 523048
rect 3292 523036 3298 523048
rect 86310 523036 86316 523048
rect 3292 523008 86316 523036
rect 3292 522996 3298 523008
rect 86310 522996 86316 523008
rect 86368 522996 86374 523048
rect 562318 522996 562324 523048
rect 562376 523036 562382 523048
rect 580166 523036 580172 523048
rect 562376 523008 580172 523036
rect 562376 522996 562382 523008
rect 580166 522996 580172 523008
rect 580224 522996 580230 523048
rect 3418 520276 3424 520328
rect 3476 520316 3482 520328
rect 121454 520316 121460 520328
rect 3476 520288 121460 520316
rect 3476 520276 3482 520288
rect 121454 520276 121460 520288
rect 121512 520276 121518 520328
rect 574830 520276 574836 520328
rect 574888 520316 574894 520328
rect 579706 520316 579712 520328
rect 574888 520288 579712 520316
rect 574888 520276 574894 520288
rect 579706 520276 579712 520288
rect 579764 520276 579770 520328
rect 3418 516128 3424 516180
rect 3476 516168 3482 516180
rect 102962 516168 102968 516180
rect 3476 516140 102968 516168
rect 3476 516128 3482 516140
rect 102962 516128 102968 516140
rect 103020 516128 103026 516180
rect 573358 516128 573364 516180
rect 573416 516168 573422 516180
rect 580166 516168 580172 516180
rect 573416 516140 580172 516168
rect 573416 516128 573422 516140
rect 580166 516128 580172 516140
rect 580224 516128 580230 516180
rect 3418 511980 3424 512032
rect 3476 512020 3482 512032
rect 96338 512020 96344 512032
rect 3476 511992 96344 512020
rect 3476 511980 3482 511992
rect 96338 511980 96344 511992
rect 96396 511980 96402 512032
rect 566550 511980 566556 512032
rect 566608 512020 566614 512032
rect 579614 512020 579620 512032
rect 566608 511992 579620 512020
rect 566608 511980 566614 511992
rect 579614 511980 579620 511992
rect 579672 511980 579678 512032
rect 3418 507832 3424 507884
rect 3476 507872 3482 507884
rect 109678 507872 109684 507884
rect 3476 507844 109684 507872
rect 3476 507832 3482 507844
rect 109678 507832 109684 507844
rect 109736 507832 109742 507884
rect 558178 507832 558184 507884
rect 558236 507872 558242 507884
rect 580166 507872 580172 507884
rect 558236 507844 580172 507872
rect 558236 507832 558242 507844
rect 580166 507832 580172 507844
rect 580224 507832 580230 507884
rect 3234 503684 3240 503736
rect 3292 503724 3298 503736
rect 120810 503724 120816 503736
rect 3292 503696 120816 503724
rect 3292 503684 3298 503696
rect 120810 503684 120816 503696
rect 120868 503684 120874 503736
rect 192570 503684 192576 503736
rect 192628 503724 192634 503736
rect 580074 503724 580080 503736
rect 192628 503696 580080 503724
rect 192628 503684 192634 503696
rect 580074 503684 580080 503696
rect 580132 503684 580138 503736
rect 3326 499536 3332 499588
rect 3384 499576 3390 499588
rect 97350 499576 97356 499588
rect 3384 499548 97356 499576
rect 3384 499536 3390 499548
rect 97350 499536 97356 499548
rect 97408 499536 97414 499588
rect 576302 499536 576308 499588
rect 576360 499576 576366 499588
rect 580166 499576 580172 499588
rect 576360 499548 580172 499576
rect 576360 499536 576366 499548
rect 580166 499536 580172 499548
rect 580224 499536 580230 499588
rect 2866 495456 2872 495508
rect 2924 495496 2930 495508
rect 93210 495496 93216 495508
rect 2924 495468 93216 495496
rect 2924 495456 2930 495468
rect 93210 495456 93216 495468
rect 93268 495456 93274 495508
rect 558270 495456 558276 495508
rect 558328 495496 558334 495508
rect 580166 495496 580172 495508
rect 558328 495468 580172 495496
rect 558328 495456 558334 495468
rect 580166 495456 580172 495468
rect 580224 495456 580230 495508
rect 3418 491308 3424 491360
rect 3476 491348 3482 491360
rect 109770 491348 109776 491360
rect 3476 491320 109776 491348
rect 3476 491308 3482 491320
rect 109770 491308 109776 491320
rect 109828 491308 109834 491360
rect 3418 487160 3424 487212
rect 3476 487200 3482 487212
rect 14458 487200 14464 487212
rect 3476 487172 14464 487200
rect 3476 487160 3482 487172
rect 14458 487160 14464 487172
rect 14516 487160 14522 487212
rect 569218 487160 569224 487212
rect 569276 487200 569282 487212
rect 580166 487200 580172 487212
rect 569276 487172 580172 487200
rect 569276 487160 569282 487172
rect 580166 487160 580172 487172
rect 580224 487160 580230 487212
rect 3510 483012 3516 483064
rect 3568 483052 3574 483064
rect 17218 483052 17224 483064
rect 3568 483024 17224 483052
rect 3568 483012 3574 483024
rect 17218 483012 17224 483024
rect 17276 483012 17282 483064
rect 182174 483012 182180 483064
rect 182232 483052 182238 483064
rect 580166 483052 580172 483064
rect 182232 483024 580172 483052
rect 182232 483012 182238 483024
rect 580166 483012 580172 483024
rect 580224 483012 580230 483064
rect 3418 478864 3424 478916
rect 3476 478904 3482 478916
rect 91830 478904 91836 478916
rect 3476 478876 91836 478904
rect 3476 478864 3482 478876
rect 91830 478864 91836 478876
rect 91888 478864 91894 478916
rect 563698 478864 563704 478916
rect 563756 478904 563762 478916
rect 580166 478904 580172 478916
rect 563756 478876 580172 478904
rect 563756 478864 563762 478876
rect 580166 478864 580172 478876
rect 580224 478864 580230 478916
rect 3234 474716 3240 474768
rect 3292 474756 3298 474768
rect 120074 474756 120080 474768
rect 3292 474728 120080 474756
rect 3292 474716 3298 474728
rect 120074 474716 120080 474728
rect 120132 474716 120138 474768
rect 561030 474716 561036 474768
rect 561088 474756 561094 474768
rect 580166 474756 580172 474768
rect 561088 474728 580172 474756
rect 561088 474716 561094 474728
rect 580166 474716 580172 474728
rect 580224 474716 580230 474768
rect 3418 471996 3424 472048
rect 3476 472036 3482 472048
rect 107194 472036 107200 472048
rect 3476 472008 107200 472036
rect 3476 471996 3482 472008
rect 107194 471996 107200 472008
rect 107252 471996 107258 472048
rect 561122 471996 561128 472048
rect 561180 472036 561186 472048
rect 580166 472036 580172 472048
rect 561180 472008 580172 472036
rect 561180 471996 561186 472008
rect 580166 471996 580172 472008
rect 580224 471996 580230 472048
rect 3418 467848 3424 467900
rect 3476 467888 3482 467900
rect 131114 467888 131120 467900
rect 3476 467860 131120 467888
rect 3476 467848 3482 467860
rect 131114 467848 131120 467860
rect 131172 467848 131178 467900
rect 563790 467848 563796 467900
rect 563848 467888 563854 467900
rect 580166 467888 580172 467900
rect 563848 467860 580172 467888
rect 563848 467848 563854 467860
rect 580166 467848 580172 467860
rect 580224 467848 580230 467900
rect 3418 463700 3424 463752
rect 3476 463740 3482 463752
rect 107102 463740 107108 463752
rect 3476 463712 107108 463740
rect 3476 463700 3482 463712
rect 107102 463700 107108 463712
rect 107160 463700 107166 463752
rect 562410 463700 562416 463752
rect 562468 463740 562474 463752
rect 580166 463740 580172 463752
rect 562468 463712 580172 463740
rect 562468 463700 562474 463712
rect 580166 463700 580172 463712
rect 580224 463700 580230 463752
rect 3418 459552 3424 459604
rect 3476 459592 3482 459604
rect 100110 459592 100116 459604
rect 3476 459564 100116 459592
rect 3476 459552 3482 459564
rect 100110 459552 100116 459564
rect 100168 459552 100174 459604
rect 552842 459552 552848 459604
rect 552900 459592 552906 459604
rect 580166 459592 580172 459604
rect 552900 459564 580172 459592
rect 552900 459552 552906 459564
rect 580166 459552 580172 459564
rect 580224 459552 580230 459604
rect 3234 455404 3240 455456
rect 3292 455444 3298 455456
rect 94682 455444 94688 455456
rect 3292 455416 94688 455444
rect 3292 455404 3298 455416
rect 94682 455404 94688 455416
rect 94740 455404 94746 455456
rect 558362 455404 558368 455456
rect 558420 455444 558426 455456
rect 580074 455444 580080 455456
rect 558420 455416 580080 455444
rect 558420 455404 558426 455416
rect 580074 455404 580080 455416
rect 580132 455404 580138 455456
rect 3326 451256 3332 451308
rect 3384 451296 3390 451308
rect 103606 451296 103612 451308
rect 3384 451268 103612 451296
rect 3384 451256 3390 451268
rect 103606 451256 103612 451268
rect 103664 451256 103670 451308
rect 124858 451256 124864 451308
rect 124916 451296 124922 451308
rect 580166 451296 580172 451308
rect 124916 451268 580172 451296
rect 124916 451256 124922 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 572070 447108 572076 447160
rect 572128 447148 572134 447160
rect 579706 447148 579712 447160
rect 572128 447120 579712 447148
rect 572128 447108 572134 447120
rect 579706 447108 579712 447120
rect 579764 447108 579770 447160
rect 3418 442960 3424 443012
rect 3476 443000 3482 443012
rect 86402 443000 86408 443012
rect 3476 442972 86408 443000
rect 3476 442960 3482 442972
rect 86402 442960 86408 442972
rect 86460 442960 86466 443012
rect 561214 442960 561220 443012
rect 561272 443000 561278 443012
rect 580166 443000 580172 443012
rect 561272 442972 580172 443000
rect 561272 442960 561278 442972
rect 580166 442960 580172 442972
rect 580224 442960 580230 443012
rect 570782 434732 570788 434784
rect 570840 434772 570846 434784
rect 580166 434772 580172 434784
rect 570840 434744 580172 434772
rect 570840 434732 570846 434744
rect 580166 434732 580172 434744
rect 580224 434732 580230 434784
rect 3510 430584 3516 430636
rect 3568 430624 3574 430636
rect 89162 430624 89168 430636
rect 3568 430596 89168 430624
rect 3568 430584 3574 430596
rect 89162 430584 89168 430596
rect 89220 430584 89226 430636
rect 568022 430584 568028 430636
rect 568080 430624 568086 430636
rect 580166 430624 580172 430636
rect 568080 430596 580172 430624
rect 568080 430584 568086 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 2866 426436 2872 426488
rect 2924 426476 2930 426488
rect 103054 426476 103060 426488
rect 2924 426448 103060 426476
rect 2924 426436 2930 426448
rect 103054 426436 103060 426448
rect 103112 426436 103118 426488
rect 563882 426436 563888 426488
rect 563940 426476 563946 426488
rect 580166 426476 580172 426488
rect 563940 426448 580172 426476
rect 563940 426436 563946 426448
rect 580166 426436 580172 426448
rect 580224 426436 580230 426488
rect 574922 423648 574928 423700
rect 574980 423688 574986 423700
rect 580166 423688 580172 423700
rect 574980 423660 580172 423688
rect 574980 423648 574986 423660
rect 580166 423648 580172 423660
rect 580224 423648 580230 423700
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 98914 422328 98920 422340
rect 3016 422300 98920 422328
rect 3016 422288 3022 422300
rect 98914 422288 98920 422300
rect 98972 422288 98978 422340
rect 3510 419500 3516 419552
rect 3568 419540 3574 419552
rect 103146 419540 103152 419552
rect 3568 419512 103152 419540
rect 3568 419500 3574 419512
rect 103146 419500 103152 419512
rect 103204 419500 103210 419552
rect 191742 419500 191748 419552
rect 191800 419540 191806 419552
rect 580166 419540 580172 419552
rect 191800 419512 580172 419540
rect 191800 419500 191806 419512
rect 580166 419500 580172 419512
rect 580224 419500 580230 419552
rect 3510 415420 3516 415472
rect 3568 415460 3574 415472
rect 108298 415460 108304 415472
rect 3568 415432 108304 415460
rect 3568 415420 3574 415432
rect 108298 415420 108304 415432
rect 108356 415420 108362 415472
rect 210418 415420 210424 415472
rect 210476 415460 210482 415472
rect 580166 415460 580172 415472
rect 210476 415432 580172 415460
rect 210476 415420 210482 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 3510 411272 3516 411324
rect 3568 411312 3574 411324
rect 90542 411312 90548 411324
rect 3568 411284 90548 411312
rect 3568 411272 3574 411284
rect 90542 411272 90548 411284
rect 90600 411272 90606 411324
rect 575106 411272 575112 411324
rect 575164 411312 575170 411324
rect 579982 411312 579988 411324
rect 575164 411284 579988 411312
rect 575164 411272 575170 411284
rect 579982 411272 579988 411284
rect 580040 411272 580046 411324
rect 3510 407124 3516 407176
rect 3568 407164 3574 407176
rect 93302 407164 93308 407176
rect 3568 407136 93308 407164
rect 3568 407124 3574 407136
rect 93302 407124 93308 407136
rect 93360 407124 93366 407176
rect 124214 407124 124220 407176
rect 124272 407164 124278 407176
rect 580166 407164 580172 407176
rect 124272 407136 580172 407164
rect 124272 407124 124278 407136
rect 580166 407124 580172 407136
rect 580224 407124 580230 407176
rect 3326 402976 3332 403028
rect 3384 403016 3390 403028
rect 96154 403016 96160 403028
rect 3384 402988 96160 403016
rect 3384 402976 3390 402988
rect 96154 402976 96160 402988
rect 96212 402976 96218 403028
rect 565170 402976 565176 403028
rect 565228 403016 565234 403028
rect 580166 403016 580172 403028
rect 565228 402988 580172 403016
rect 565228 402976 565234 402988
rect 580166 402976 580172 402988
rect 580224 402976 580230 403028
rect 179414 398828 179420 398880
rect 179472 398868 179478 398880
rect 579706 398868 579712 398880
rect 179472 398840 579712 398868
rect 179472 398828 179478 398840
rect 579706 398828 579712 398840
rect 579764 398828 579770 398880
rect 576394 394680 576400 394732
rect 576452 394720 576458 394732
rect 580166 394720 580172 394732
rect 576452 394692 580172 394720
rect 576452 394680 576458 394692
rect 580166 394680 580172 394692
rect 580224 394680 580230 394732
rect 3510 390532 3516 390584
rect 3568 390572 3574 390584
rect 118694 390572 118700 390584
rect 3568 390544 118700 390572
rect 3568 390532 3574 390544
rect 118694 390532 118700 390544
rect 118752 390532 118758 390584
rect 572162 390532 572168 390584
rect 572220 390572 572226 390584
rect 580166 390572 580172 390584
rect 572220 390544 580172 390572
rect 572220 390532 572226 390544
rect 580166 390532 580172 390544
rect 580224 390532 580230 390584
rect 3510 386384 3516 386436
rect 3568 386424 3574 386436
rect 100202 386424 100208 386436
rect 3568 386396 100208 386424
rect 3568 386384 3574 386396
rect 100202 386384 100208 386396
rect 100260 386384 100266 386436
rect 189810 386384 189816 386436
rect 189868 386424 189874 386436
rect 580166 386424 580172 386436
rect 189868 386396 580172 386424
rect 189868 386384 189874 386396
rect 580166 386384 580172 386396
rect 580224 386384 580230 386436
rect 2866 378156 2872 378208
rect 2924 378196 2930 378208
rect 89254 378196 89260 378208
rect 2924 378168 89260 378196
rect 2924 378156 2930 378168
rect 89254 378156 89260 378168
rect 89312 378156 89318 378208
rect 184934 375368 184940 375420
rect 184992 375408 184998 375420
rect 580166 375408 580172 375420
rect 184992 375380 580172 375408
rect 184992 375368 184998 375380
rect 580166 375368 580172 375380
rect 580224 375368 580230 375420
rect 2958 374008 2964 374060
rect 3016 374048 3022 374060
rect 108390 374048 108396 374060
rect 3016 374020 108396 374048
rect 3016 374008 3022 374020
rect 108390 374008 108396 374020
rect 108448 374008 108454 374060
rect 555418 371220 555424 371272
rect 555476 371260 555482 371272
rect 579798 371260 579804 371272
rect 555476 371232 579804 371260
rect 555476 371220 555482 371232
rect 579798 371220 579804 371232
rect 579856 371220 579862 371272
rect 3050 369860 3056 369912
rect 3108 369900 3114 369912
rect 111150 369900 111156 369912
rect 3108 369872 111156 369900
rect 3108 369860 3114 369872
rect 111150 369860 111156 369872
rect 111208 369860 111214 369912
rect 189902 367072 189908 367124
rect 189960 367112 189966 367124
rect 580166 367112 580172 367124
rect 189960 367084 580172 367112
rect 189960 367072 189966 367084
rect 580166 367072 580172 367084
rect 580224 367072 580230 367124
rect 3050 361564 3056 361616
rect 3108 361604 3114 361616
rect 97442 361604 97448 361616
rect 3108 361576 97448 361604
rect 3108 361564 3114 361576
rect 97442 361564 97448 361576
rect 97500 361564 97506 361616
rect 3326 358776 3332 358828
rect 3384 358816 3390 358828
rect 105630 358816 105636 358828
rect 3384 358788 105636 358816
rect 3384 358776 3390 358788
rect 105630 358776 105636 358788
rect 105688 358776 105694 358828
rect 566734 358776 566740 358828
rect 566792 358816 566798 358828
rect 580166 358816 580172 358828
rect 566792 358788 580172 358816
rect 566792 358776 566798 358788
rect 580166 358776 580172 358788
rect 580224 358776 580230 358828
rect 3326 354696 3332 354748
rect 3384 354736 3390 354748
rect 100294 354736 100300 354748
rect 3384 354708 100300 354736
rect 3384 354696 3390 354708
rect 100294 354696 100300 354708
rect 100352 354696 100358 354748
rect 178034 354696 178040 354748
rect 178092 354736 178098 354748
rect 580166 354736 580172 354748
rect 178092 354708 580172 354736
rect 178092 354696 178098 354708
rect 580166 354696 580172 354708
rect 580224 354696 580230 354748
rect 3510 350548 3516 350600
rect 3568 350588 3574 350600
rect 104250 350588 104256 350600
rect 3568 350560 104256 350588
rect 3568 350548 3574 350560
rect 104250 350548 104256 350560
rect 104308 350548 104314 350600
rect 206278 350548 206284 350600
rect 206336 350588 206342 350600
rect 580166 350588 580172 350600
rect 206336 350560 580172 350588
rect 206336 350548 206342 350560
rect 580166 350548 580172 350560
rect 580224 350548 580230 350600
rect 3326 346400 3332 346452
rect 3384 346440 3390 346452
rect 75178 346440 75184 346452
rect 3384 346412 75184 346440
rect 3384 346400 3390 346412
rect 75178 346400 75184 346412
rect 75236 346400 75242 346452
rect 569310 346400 569316 346452
rect 569368 346440 569374 346452
rect 580166 346440 580172 346452
rect 569368 346412 580172 346440
rect 569368 346400 569374 346412
rect 580166 346400 580172 346412
rect 580224 346400 580230 346452
rect 3510 342252 3516 342304
rect 3568 342292 3574 342304
rect 104894 342292 104900 342304
rect 3568 342264 104900 342292
rect 3568 342252 3574 342264
rect 104894 342252 104900 342264
rect 104952 342252 104958 342304
rect 563974 342252 563980 342304
rect 564032 342292 564038 342304
rect 579706 342292 579712 342304
rect 564032 342264 579712 342292
rect 564032 342252 564038 342264
rect 579706 342252 579712 342264
rect 579764 342252 579770 342304
rect 3510 338104 3516 338156
rect 3568 338144 3574 338156
rect 108482 338144 108488 338156
rect 3568 338116 108488 338144
rect 3568 338104 3574 338116
rect 108482 338104 108488 338116
rect 108540 338104 108546 338156
rect 577590 338104 577596 338156
rect 577648 338144 577654 338156
rect 579614 338144 579620 338156
rect 577648 338116 579620 338144
rect 577648 338104 577654 338116
rect 579614 338104 579620 338116
rect 579672 338104 579678 338156
rect 572254 331236 572260 331288
rect 572312 331276 572318 331288
rect 579706 331276 579712 331288
rect 572312 331248 579712 331276
rect 572312 331236 572318 331248
rect 579706 331236 579712 331248
rect 579764 331236 579770 331288
rect 2958 329808 2964 329860
rect 3016 329848 3022 329860
rect 109862 329848 109868 329860
rect 3016 329820 109868 329848
rect 3016 329808 3022 329820
rect 109862 329808 109868 329820
rect 109920 329808 109926 329860
rect 3050 321580 3056 321632
rect 3108 321620 3114 321632
rect 94774 321620 94780 321632
rect 3108 321592 94780 321620
rect 3108 321580 3114 321592
rect 94774 321580 94780 321592
rect 94832 321580 94838 321632
rect 577682 318792 577688 318844
rect 577740 318832 577746 318844
rect 579706 318832 579712 318844
rect 577740 318804 579712 318832
rect 577740 318792 577746 318804
rect 579706 318792 579712 318804
rect 579764 318792 579770 318844
rect 3510 317432 3516 317484
rect 3568 317472 3574 317484
rect 94866 317472 94872 317484
rect 3568 317444 94872 317472
rect 3568 317432 3574 317444
rect 94866 317432 94872 317444
rect 94924 317432 94930 317484
rect 575014 314644 575020 314696
rect 575072 314684 575078 314696
rect 579614 314684 579620 314696
rect 575072 314656 579620 314684
rect 575072 314644 575078 314656
rect 579614 314644 579620 314656
rect 579672 314644 579678 314696
rect 3050 313284 3056 313336
rect 3108 313324 3114 313336
rect 126974 313324 126980 313336
rect 3108 313296 126980 313324
rect 3108 313284 3114 313296
rect 126974 313284 126980 313296
rect 127032 313284 127038 313336
rect 558454 310496 558460 310548
rect 558512 310536 558518 310548
rect 580166 310536 580172 310548
rect 558512 310508 580172 310536
rect 558512 310496 558518 310508
rect 580166 310496 580172 310508
rect 580224 310496 580230 310548
rect 3142 309136 3148 309188
rect 3200 309176 3206 309188
rect 108574 309176 108580 309188
rect 3200 309148 108580 309176
rect 3200 309136 3206 309148
rect 108574 309136 108580 309148
rect 108632 309136 108638 309188
rect 564066 306348 564072 306400
rect 564124 306388 564130 306400
rect 580166 306388 580172 306400
rect 564124 306360 580172 306388
rect 564124 306348 564130 306360
rect 580166 306348 580172 306360
rect 580224 306348 580230 306400
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 105722 305028 105728 305040
rect 3292 305000 105728 305028
rect 3292 304988 3298 305000
rect 105722 304988 105728 305000
rect 105780 304988 105786 305040
rect 569402 302200 569408 302252
rect 569460 302240 569466 302252
rect 580166 302240 580172 302252
rect 569460 302212 580172 302240
rect 569460 302200 569466 302212
rect 580166 302200 580172 302212
rect 580224 302200 580230 302252
rect 3142 300840 3148 300892
rect 3200 300880 3206 300892
rect 118786 300880 118792 300892
rect 3200 300852 118792 300880
rect 3200 300840 3206 300852
rect 118786 300840 118792 300852
rect 118844 300840 118850 300892
rect 3326 298120 3332 298172
rect 3384 298160 3390 298172
rect 118050 298160 118056 298172
rect 3384 298132 118056 298160
rect 3384 298120 3390 298132
rect 118050 298120 118056 298132
rect 118108 298120 118114 298172
rect 3510 293972 3516 294024
rect 3568 294012 3574 294024
rect 101490 294012 101496 294024
rect 3568 293984 101496 294012
rect 3568 293972 3574 293984
rect 101490 293972 101496 293984
rect 101548 293972 101554 294024
rect 170398 293972 170404 294024
rect 170456 294012 170462 294024
rect 580166 294012 580172 294024
rect 170456 293984 580172 294012
rect 170456 293972 170462 293984
rect 580166 293972 580172 293984
rect 580224 293972 580230 294024
rect 3510 289824 3516 289876
rect 3568 289864 3574 289876
rect 120258 289864 120264 289876
rect 3568 289836 120264 289864
rect 3568 289824 3574 289836
rect 120258 289824 120264 289836
rect 120316 289824 120322 289876
rect 558546 289824 558552 289876
rect 558604 289864 558610 289876
rect 579982 289864 579988 289876
rect 558604 289836 579988 289864
rect 558604 289824 558610 289836
rect 579982 289824 579988 289836
rect 580040 289824 580046 289876
rect 2866 285676 2872 285728
rect 2924 285716 2930 285728
rect 108666 285716 108672 285728
rect 2924 285688 108672 285716
rect 2924 285676 2930 285688
rect 108666 285676 108672 285688
rect 108724 285676 108730 285728
rect 572346 285676 572352 285728
rect 572404 285716 572410 285728
rect 579982 285716 579988 285728
rect 572404 285688 579988 285716
rect 572404 285676 572410 285688
rect 579982 285676 579988 285688
rect 580040 285676 580046 285728
rect 555510 282888 555516 282940
rect 555568 282928 555574 282940
rect 580166 282928 580172 282940
rect 555568 282900 580172 282928
rect 555568 282888 555574 282900
rect 580166 282888 580172 282900
rect 580224 282888 580230 282940
rect 2958 281528 2964 281580
rect 3016 281568 3022 281580
rect 102686 281568 102692 281580
rect 3016 281540 102692 281568
rect 3016 281528 3022 281540
rect 102686 281528 102692 281540
rect 102744 281528 102750 281580
rect 561306 278740 561312 278792
rect 561364 278780 561370 278792
rect 580166 278780 580172 278792
rect 561364 278752 580172 278780
rect 561364 278740 561370 278752
rect 580166 278740 580172 278752
rect 580224 278740 580230 278792
rect 122926 277992 122932 278044
rect 122984 278032 122990 278044
rect 498838 278032 498844 278044
rect 122984 278004 498844 278032
rect 122984 277992 122990 278004
rect 498838 277992 498844 278004
rect 498896 277992 498902 278044
rect 3050 277380 3056 277432
rect 3108 277420 3114 277432
rect 97810 277420 97816 277432
rect 3108 277392 97816 277420
rect 3108 277380 3114 277392
rect 97810 277380 97816 277392
rect 97868 277380 97874 277432
rect 195238 276632 195244 276684
rect 195296 276672 195302 276684
rect 524414 276672 524420 276684
rect 195296 276644 524420 276672
rect 195296 276632 195302 276644
rect 524414 276632 524420 276644
rect 524472 276632 524478 276684
rect 169754 276020 169760 276072
rect 169812 276060 169818 276072
rect 195238 276060 195244 276072
rect 169812 276032 195244 276060
rect 169812 276020 169818 276032
rect 195238 276020 195244 276032
rect 195296 276020 195302 276072
rect 566826 274660 566832 274712
rect 566884 274700 566890 274712
rect 580166 274700 580172 274712
rect 566884 274672 580172 274700
rect 566884 274660 566890 274672
rect 580166 274660 580172 274672
rect 580224 274660 580230 274712
rect 147674 273912 147680 273964
rect 147732 273952 147738 273964
rect 218054 273952 218060 273964
rect 147732 273924 218060 273952
rect 147732 273912 147738 273924
rect 218054 273912 218060 273924
rect 218112 273912 218118 273964
rect 3510 273232 3516 273284
rect 3568 273272 3574 273284
rect 99926 273272 99932 273284
rect 3568 273244 99932 273272
rect 3568 273232 3574 273244
rect 99926 273232 99932 273244
rect 99984 273232 99990 273284
rect 191650 272484 191656 272536
rect 191708 272524 191714 272536
rect 206278 272524 206284 272536
rect 191708 272496 206284 272524
rect 191708 272484 191714 272496
rect 206278 272484 206284 272496
rect 206336 272484 206342 272536
rect 155954 271872 155960 271924
rect 156012 271912 156018 271924
rect 190454 271912 190460 271924
rect 156012 271884 190460 271912
rect 156012 271872 156018 271884
rect 190454 271872 190460 271884
rect 190512 271912 190518 271924
rect 191650 271912 191656 271924
rect 190512 271884 191656 271912
rect 190512 271872 190518 271884
rect 191650 271872 191656 271884
rect 191708 271872 191714 271924
rect 149146 271192 149152 271244
rect 149204 271232 149210 271244
rect 202138 271232 202144 271244
rect 149204 271204 202144 271232
rect 149204 271192 149210 271204
rect 202138 271192 202144 271204
rect 202196 271192 202202 271244
rect 17218 271124 17224 271176
rect 17276 271164 17282 271176
rect 110506 271164 110512 271176
rect 17276 271136 110512 271164
rect 17276 271124 17282 271136
rect 110506 271124 110512 271136
rect 110564 271124 110570 271176
rect 142798 271124 142804 271176
rect 142856 271164 142862 271176
rect 230474 271164 230480 271176
rect 142856 271136 230480 271164
rect 142856 271124 142862 271136
rect 230474 271124 230480 271136
rect 230532 271124 230538 271176
rect 110506 270512 110512 270564
rect 110564 270552 110570 270564
rect 111702 270552 111708 270564
rect 110564 270524 111708 270552
rect 110564 270512 110570 270524
rect 111702 270512 111708 270524
rect 111760 270552 111766 270564
rect 133966 270552 133972 270564
rect 111760 270524 133972 270552
rect 111760 270512 111766 270524
rect 133966 270512 133972 270524
rect 134024 270512 134030 270564
rect 577866 270512 577872 270564
rect 577924 270552 577930 270564
rect 579706 270552 579712 270564
rect 577924 270524 579712 270552
rect 577924 270512 577930 270524
rect 579706 270512 579712 270524
rect 579764 270512 579770 270564
rect 132586 269764 132592 269816
rect 132644 269804 132650 269816
rect 200758 269804 200764 269816
rect 132644 269776 200764 269804
rect 132644 269764 132650 269776
rect 200758 269764 200764 269776
rect 200816 269764 200822 269816
rect 3050 269084 3056 269136
rect 3108 269124 3114 269136
rect 183646 269124 183652 269136
rect 3108 269096 183652 269124
rect 3108 269084 3114 269096
rect 183646 269084 183652 269096
rect 183704 269084 183710 269136
rect 10318 268404 10324 268456
rect 10376 268444 10382 268456
rect 160094 268444 160100 268456
rect 10376 268416 160100 268444
rect 10376 268404 10382 268416
rect 160094 268404 160100 268416
rect 160152 268404 160158 268456
rect 145006 268336 145012 268388
rect 145064 268376 145070 268388
rect 472618 268376 472624 268388
rect 145064 268348 472624 268376
rect 145064 268336 145070 268348
rect 472618 268336 472624 268348
rect 472676 268336 472682 268388
rect 111058 267724 111064 267776
rect 111116 267764 111122 267776
rect 114462 267764 114468 267776
rect 111116 267736 114468 267764
rect 111116 267724 111122 267736
rect 114462 267724 114468 267736
rect 114520 267764 114526 267776
rect 139486 267764 139492 267776
rect 114520 267736 139492 267764
rect 114520 267724 114526 267736
rect 139486 267724 139492 267736
rect 139544 267724 139550 267776
rect 144822 267044 144828 267096
rect 144880 267084 144886 267096
rect 170398 267084 170404 267096
rect 144880 267056 170404 267084
rect 144880 267044 144886 267056
rect 170398 267044 170404 267056
rect 170456 267044 170462 267096
rect 7558 266976 7564 267028
rect 7616 267016 7622 267028
rect 167454 267016 167460 267028
rect 7616 266988 167460 267016
rect 7616 266976 7622 266988
rect 167454 266976 167460 266988
rect 167512 266976 167518 267028
rect 196986 266636 196992 266688
rect 197044 266676 197050 266688
rect 197998 266676 198004 266688
rect 197044 266648 198004 266676
rect 197044 266636 197050 266648
rect 197998 266636 198004 266648
rect 198056 266636 198062 266688
rect 169754 266432 169760 266484
rect 169812 266472 169818 266484
rect 198734 266472 198740 266484
rect 169812 266444 198740 266472
rect 169812 266432 169818 266444
rect 198734 266432 198740 266444
rect 198792 266472 198798 266484
rect 198792 266444 200114 266472
rect 198792 266432 198798 266444
rect 163958 266364 163964 266416
rect 164016 266404 164022 266416
rect 196986 266404 196992 266416
rect 164016 266376 196992 266404
rect 164016 266364 164022 266376
rect 196986 266364 196992 266376
rect 197044 266364 197050 266416
rect 200086 266404 200114 266444
rect 579614 266404 579620 266416
rect 200086 266376 579620 266404
rect 579614 266364 579620 266376
rect 579672 266364 579678 266416
rect 189074 265956 189080 266008
rect 189132 265996 189138 266008
rect 210418 265996 210424 266008
rect 189132 265968 210424 265996
rect 189132 265956 189138 265968
rect 210418 265956 210424 265968
rect 210476 265956 210482 266008
rect 161474 265888 161480 265940
rect 161532 265928 161538 265940
rect 189994 265928 190000 265940
rect 161532 265900 190000 265928
rect 161532 265888 161538 265900
rect 189994 265888 190000 265900
rect 190052 265888 190058 265940
rect 153194 265820 153200 265872
rect 153252 265860 153258 265872
rect 197354 265860 197360 265872
rect 153252 265832 197360 265860
rect 153252 265820 153258 265832
rect 197354 265820 197360 265832
rect 197412 265820 197418 265872
rect 133874 265752 133880 265804
rect 133932 265792 133938 265804
rect 189626 265792 189632 265804
rect 133932 265764 189632 265792
rect 133932 265752 133938 265764
rect 189626 265752 189632 265764
rect 189684 265752 189690 265804
rect 136542 265684 136548 265736
rect 136600 265724 136606 265736
rect 193858 265724 193864 265736
rect 136600 265696 193864 265724
rect 136600 265684 136606 265696
rect 193858 265684 193864 265696
rect 193916 265684 193922 265736
rect 148042 265616 148048 265668
rect 148100 265656 148106 265668
rect 492674 265656 492680 265668
rect 148100 265628 492680 265656
rect 148100 265616 148106 265628
rect 492674 265616 492680 265628
rect 492732 265616 492738 265668
rect 3142 264936 3148 264988
rect 3200 264976 3206 264988
rect 106826 264976 106832 264988
rect 3200 264948 106832 264976
rect 3200 264936 3206 264948
rect 106826 264936 106832 264948
rect 106884 264936 106890 264988
rect 118142 264936 118148 264988
rect 118200 264976 118206 264988
rect 151906 264976 151912 264988
rect 118200 264948 151912 264976
rect 118200 264936 118206 264948
rect 151906 264936 151912 264948
rect 151964 264936 151970 264988
rect 154482 264936 154488 264988
rect 154540 264976 154546 264988
rect 189074 264976 189080 264988
rect 154540 264948 189080 264976
rect 154540 264936 154546 264948
rect 189074 264936 189080 264948
rect 189132 264976 189138 264988
rect 189534 264976 189540 264988
rect 189132 264948 189540 264976
rect 189132 264936 189138 264948
rect 189534 264936 189540 264948
rect 189592 264936 189598 264988
rect 146202 264392 146208 264444
rect 146260 264432 146266 264444
rect 192570 264432 192576 264444
rect 146260 264404 192576 264432
rect 146260 264392 146266 264404
rect 192570 264392 192576 264404
rect 192628 264392 192634 264444
rect 75178 264324 75184 264376
rect 75236 264364 75242 264376
rect 158714 264364 158720 264376
rect 75236 264336 158720 264364
rect 75236 264324 75242 264336
rect 158714 264324 158720 264336
rect 158772 264324 158778 264376
rect 14458 264256 14464 264308
rect 14516 264296 14522 264308
rect 158346 264296 158352 264308
rect 14516 264268 158352 264296
rect 14516 264256 14522 264268
rect 158346 264256 158352 264268
rect 158404 264256 158410 264308
rect 149238 264188 149244 264240
rect 149296 264228 149302 264240
rect 150342 264228 150348 264240
rect 149296 264200 150348 264228
rect 149296 264188 149302 264200
rect 150342 264188 150348 264200
rect 150400 264228 150406 264240
rect 400858 264228 400864 264240
rect 150400 264200 400864 264228
rect 150400 264188 150406 264200
rect 400858 264188 400864 264200
rect 400916 264188 400922 264240
rect 115750 263984 115756 264036
rect 115808 264024 115814 264036
rect 124858 264024 124864 264036
rect 115808 263996 124864 264024
rect 115808 263984 115814 263996
rect 124858 263984 124864 263996
rect 124916 264024 124922 264036
rect 125226 264024 125232 264036
rect 124916 263996 125232 264024
rect 124916 263984 124922 263996
rect 125226 263984 125232 263996
rect 125284 263984 125290 264036
rect 117130 263916 117136 263968
rect 117188 263956 117194 263968
rect 126974 263956 126980 263968
rect 117188 263928 126980 263956
rect 117188 263916 117194 263928
rect 126974 263916 126980 263928
rect 127032 263956 127038 263968
rect 127710 263956 127716 263968
rect 127032 263928 127716 263956
rect 127032 263916 127038 263928
rect 127710 263916 127716 263928
rect 127768 263916 127774 263968
rect 114186 263848 114192 263900
rect 114244 263888 114250 263900
rect 132586 263888 132592 263900
rect 114244 263860 132592 263888
rect 114244 263848 114250 263860
rect 132586 263848 132592 263860
rect 132644 263888 132650 263900
rect 133506 263888 133512 263900
rect 132644 263860 133512 263888
rect 132644 263848 132650 263860
rect 133506 263848 133512 263860
rect 133564 263848 133570 263900
rect 118510 263780 118516 263832
rect 118568 263820 118574 263832
rect 145374 263820 145380 263832
rect 118568 263792 145380 263820
rect 118568 263780 118574 263792
rect 145374 263780 145380 263792
rect 145432 263820 145438 263832
rect 146202 263820 146208 263832
rect 145432 263792 146208 263820
rect 145432 263780 145438 263792
rect 146202 263780 146208 263792
rect 146260 263780 146266 263832
rect 115658 263712 115664 263764
rect 115716 263752 115722 263764
rect 142614 263752 142620 263764
rect 115716 263724 142620 263752
rect 115716 263712 115722 263724
rect 142614 263712 142620 263724
rect 142672 263712 142678 263764
rect 166718 263712 166724 263764
rect 166776 263752 166782 263764
rect 166776 263724 180794 263752
rect 166776 263712 166782 263724
rect 119982 263644 119988 263696
rect 120040 263684 120046 263696
rect 149238 263684 149244 263696
rect 120040 263656 149244 263684
rect 120040 263644 120046 263656
rect 149238 263644 149244 263656
rect 149296 263644 149302 263696
rect 180766 263684 180794 263724
rect 198918 263684 198924 263696
rect 180766 263656 198924 263684
rect 198918 263644 198924 263656
rect 198976 263644 198982 263696
rect 112898 263576 112904 263628
rect 112956 263616 112962 263628
rect 143718 263616 143724 263628
rect 112956 263588 143724 263616
rect 112956 263576 112962 263588
rect 143718 263576 143724 263588
rect 143776 263616 143782 263628
rect 144822 263616 144828 263628
rect 143776 263588 144828 263616
rect 143776 263576 143782 263588
rect 144822 263576 144828 263588
rect 144880 263576 144886 263628
rect 158714 263576 158720 263628
rect 158772 263616 158778 263628
rect 159450 263616 159456 263628
rect 158772 263588 159456 263616
rect 158772 263576 158778 263588
rect 159450 263576 159456 263588
rect 159508 263616 159514 263628
rect 193582 263616 193588 263628
rect 159508 263588 193588 263616
rect 159508 263576 159514 263588
rect 193582 263576 193588 263588
rect 193640 263576 193646 263628
rect 132126 263508 132132 263560
rect 132184 263548 132190 263560
rect 470594 263548 470600 263560
rect 132184 263520 470600 263548
rect 132184 263508 132190 263520
rect 470594 263508 470600 263520
rect 470652 263508 470658 263560
rect 23474 263440 23480 263492
rect 23532 263480 23538 263492
rect 166718 263480 166724 263492
rect 23532 263452 166724 263480
rect 23532 263440 23538 263452
rect 166718 263440 166724 263452
rect 166776 263440 166782 263492
rect 57974 263372 57980 263424
rect 58032 263412 58038 263424
rect 161934 263412 161940 263424
rect 58032 263384 161940 263412
rect 58032 263372 58038 263384
rect 161934 263372 161940 263384
rect 161992 263372 161998 263424
rect 69014 263304 69020 263356
rect 69072 263344 69078 263356
rect 171594 263344 171600 263356
rect 69072 263316 171600 263344
rect 69072 263304 69078 263316
rect 171594 263304 171600 263316
rect 171652 263304 171658 263356
rect 157242 263100 157248 263152
rect 157300 263140 157306 263152
rect 190822 263140 190828 263152
rect 157300 263112 190828 263140
rect 157300 263100 157306 263112
rect 190822 263100 190828 263112
rect 190880 263140 190886 263152
rect 267734 263140 267740 263152
rect 190880 263112 267740 263140
rect 190880 263100 190886 263112
rect 267734 263100 267740 263112
rect 267792 263100 267798 263152
rect 130010 263032 130016 263084
rect 130068 263072 130074 263084
rect 276014 263072 276020 263084
rect 130068 263044 276020 263072
rect 130068 263032 130074 263044
rect 276014 263032 276020 263044
rect 276072 263032 276078 263084
rect 196250 262964 196256 263016
rect 196308 263004 196314 263016
rect 347774 263004 347780 263016
rect 196308 262976 347780 263004
rect 196308 262964 196314 262976
rect 347774 262964 347780 262976
rect 347832 262964 347838 263016
rect 111058 262896 111064 262948
rect 111116 262936 111122 262948
rect 126974 262936 126980 262948
rect 111116 262908 126980 262936
rect 111116 262896 111122 262908
rect 126974 262896 126980 262908
rect 127032 262896 127038 262948
rect 140774 262896 140780 262948
rect 140832 262936 140838 262948
rect 299474 262936 299480 262948
rect 140832 262908 299480 262936
rect 140832 262896 140838 262908
rect 299474 262896 299480 262908
rect 299532 262896 299538 262948
rect 121546 262828 121552 262880
rect 121604 262868 121610 262880
rect 138474 262868 138480 262880
rect 121604 262840 138480 262868
rect 121604 262828 121610 262840
rect 138474 262828 138480 262840
rect 138532 262828 138538 262880
rect 164786 262828 164792 262880
rect 164844 262868 164850 262880
rect 194594 262868 194600 262880
rect 164844 262840 194600 262868
rect 164844 262828 164850 262840
rect 194594 262828 194600 262840
rect 194652 262868 194658 262880
rect 197630 262868 197636 262880
rect 194652 262840 197636 262868
rect 194652 262828 194658 262840
rect 197630 262828 197636 262840
rect 197688 262828 197694 262880
rect 477494 262868 477500 262880
rect 200086 262840 477500 262868
rect 119798 262760 119804 262812
rect 119856 262800 119862 262812
rect 152550 262800 152556 262812
rect 119856 262772 152556 262800
rect 119856 262760 119862 262772
rect 152550 262760 152556 262772
rect 152608 262760 152614 262812
rect 155678 262760 155684 262812
rect 155736 262800 155742 262812
rect 190638 262800 190644 262812
rect 155736 262772 190644 262800
rect 155736 262760 155742 262772
rect 190638 262760 190644 262772
rect 190696 262760 190702 262812
rect 119614 262692 119620 262744
rect 119672 262732 119678 262744
rect 153378 262732 153384 262744
rect 119672 262704 153384 262732
rect 119672 262692 119678 262704
rect 153378 262692 153384 262704
rect 153436 262692 153442 262744
rect 170582 262692 170588 262744
rect 170640 262732 170646 262744
rect 191098 262732 191104 262744
rect 170640 262704 191104 262732
rect 170640 262692 170646 262704
rect 191098 262692 191104 262704
rect 191156 262692 191162 262744
rect 119890 262624 119896 262676
rect 119948 262664 119954 262676
rect 137646 262664 137652 262676
rect 119948 262636 137652 262664
rect 119948 262624 119954 262636
rect 137646 262624 137652 262636
rect 137704 262624 137710 262676
rect 174722 262624 174728 262676
rect 174780 262664 174786 262676
rect 197538 262664 197544 262676
rect 174780 262636 197544 262664
rect 174780 262624 174786 262636
rect 197538 262624 197544 262636
rect 197596 262624 197602 262676
rect 116302 262556 116308 262608
rect 116360 262596 116366 262608
rect 140130 262596 140136 262608
rect 116360 262568 140136 262596
rect 116360 262556 116366 262568
rect 140130 262556 140136 262568
rect 140188 262556 140194 262608
rect 173802 262556 173808 262608
rect 173860 262596 173866 262608
rect 199102 262596 199108 262608
rect 173860 262568 199108 262596
rect 173860 262556 173866 262568
rect 199102 262556 199108 262568
rect 199160 262596 199166 262608
rect 200086 262596 200114 262840
rect 477494 262828 477500 262840
rect 477552 262828 477558 262880
rect 199160 262568 200114 262596
rect 199160 262556 199166 262568
rect 112990 262488 112996 262540
rect 113048 262528 113054 262540
rect 136818 262528 136824 262540
rect 113048 262500 136824 262528
rect 113048 262488 113054 262500
rect 136818 262488 136824 262500
rect 136876 262488 136882 262540
rect 165522 262488 165528 262540
rect 165580 262528 165586 262540
rect 192846 262528 192852 262540
rect 165580 262500 192852 262528
rect 165580 262488 165586 262500
rect 192846 262488 192852 262500
rect 192904 262488 192910 262540
rect 115566 262420 115572 262472
rect 115624 262460 115630 262472
rect 141786 262460 141792 262472
rect 115624 262432 141792 262460
rect 115624 262420 115630 262432
rect 141786 262420 141792 262432
rect 141844 262420 141850 262472
rect 160646 262420 160652 262472
rect 160704 262460 160710 262472
rect 193306 262460 193312 262472
rect 160704 262432 193312 262460
rect 160704 262420 160710 262432
rect 193306 262420 193312 262432
rect 193364 262420 193370 262472
rect 114278 262352 114284 262404
rect 114336 262392 114342 262404
rect 140774 262392 140780 262404
rect 114336 262364 140780 262392
rect 114336 262352 114342 262364
rect 140774 262352 140780 262364
rect 140832 262352 140838 262404
rect 158162 262352 158168 262404
rect 158220 262392 158226 262404
rect 190730 262392 190736 262404
rect 158220 262364 190736 262392
rect 158220 262352 158226 262364
rect 190730 262352 190736 262364
rect 190788 262352 190794 262404
rect 118234 262284 118240 262336
rect 118292 262324 118298 262336
rect 130194 262324 130200 262336
rect 118292 262296 130200 262324
rect 118292 262284 118298 262296
rect 130194 262284 130200 262296
rect 130252 262284 130258 262336
rect 177942 262284 177948 262336
rect 178000 262324 178006 262336
rect 179414 262324 179420 262336
rect 178000 262296 179420 262324
rect 178000 262284 178006 262296
rect 179414 262284 179420 262296
rect 179472 262284 179478 262336
rect 181346 262284 181352 262336
rect 181404 262324 181410 262336
rect 196250 262324 196256 262336
rect 181404 262296 196256 262324
rect 181404 262284 181410 262296
rect 196250 262284 196256 262296
rect 196308 262284 196314 262336
rect 134886 262216 134892 262268
rect 134944 262256 134950 262268
rect 135990 262256 135996 262268
rect 134944 262228 135996 262256
rect 134944 262216 134950 262228
rect 135990 262216 135996 262228
rect 136048 262216 136054 262268
rect 173066 262216 173072 262268
rect 173124 262256 173130 262268
rect 193398 262256 193404 262268
rect 173124 262228 193404 262256
rect 173124 262216 173130 262228
rect 193398 262216 193404 262228
rect 193456 262216 193462 262268
rect 577774 262216 577780 262268
rect 577832 262256 577838 262268
rect 580258 262256 580264 262268
rect 577832 262228 580264 262256
rect 577832 262216 577838 262228
rect 580258 262216 580264 262228
rect 580316 262216 580322 262268
rect 162762 260992 162768 261044
rect 162820 261032 162826 261044
rect 162820 261004 193536 261032
rect 162820 260992 162826 261004
rect 3050 260924 3056 260976
rect 3108 260964 3114 260976
rect 109954 260964 109960 260976
rect 3108 260936 109960 260964
rect 3108 260924 3114 260936
rect 109954 260924 109960 260936
rect 110012 260924 110018 260976
rect 111334 260924 111340 260976
rect 111392 260964 111398 260976
rect 144822 260964 144828 260976
rect 111392 260936 144828 260964
rect 111392 260924 111398 260936
rect 144822 260924 144828 260936
rect 144880 260964 144886 260976
rect 192570 260964 192576 260976
rect 144880 260936 192576 260964
rect 144880 260924 144886 260936
rect 192570 260924 192576 260936
rect 192628 260924 192634 260976
rect 193508 260908 193536 261004
rect 7558 260856 7564 260908
rect 7616 260896 7622 260908
rect 176654 260896 176660 260908
rect 7616 260868 176660 260896
rect 7616 260856 7622 260868
rect 176654 260856 176660 260868
rect 176712 260896 176718 260908
rect 192386 260896 192392 260908
rect 176712 260868 192392 260896
rect 176712 260856 176718 260868
rect 192386 260856 192392 260868
rect 192444 260856 192450 260908
rect 193490 260856 193496 260908
rect 193548 260896 193554 260908
rect 498838 260896 498844 260908
rect 193548 260868 498844 260896
rect 193548 260856 193554 260868
rect 498838 260856 498844 260868
rect 498896 260856 498902 260908
rect 118418 260788 118424 260840
rect 118476 260828 118482 260840
rect 122834 260828 122840 260840
rect 118476 260800 122840 260828
rect 118476 260788 118482 260800
rect 122834 260788 122840 260800
rect 122892 260788 122898 260840
rect 129734 260788 129740 260840
rect 129792 260828 129798 260840
rect 129918 260828 129924 260840
rect 129792 260800 129924 260828
rect 129792 260788 129798 260800
rect 129918 260788 129924 260800
rect 129976 260828 129982 260840
rect 132678 260828 132684 260840
rect 129976 260800 132684 260828
rect 129976 260788 129982 260800
rect 132678 260788 132684 260800
rect 132736 260788 132742 260840
rect 161198 260312 161204 260364
rect 161256 260352 161262 260364
rect 194962 260352 194968 260364
rect 161256 260324 194968 260352
rect 161256 260312 161262 260324
rect 194962 260312 194968 260324
rect 195020 260312 195026 260364
rect 113818 260244 113824 260296
rect 113876 260284 113882 260296
rect 124398 260284 124404 260296
rect 113876 260256 124404 260284
rect 113876 260244 113882 260256
rect 124398 260244 124404 260256
rect 124456 260244 124462 260296
rect 158346 260244 158352 260296
rect 158404 260284 158410 260296
rect 193766 260284 193772 260296
rect 158404 260256 193772 260284
rect 158404 260244 158410 260256
rect 193766 260244 193772 260256
rect 193824 260244 193830 260296
rect 119706 260176 119712 260228
rect 119764 260216 119770 260228
rect 144914 260216 144920 260228
rect 119764 260188 144920 260216
rect 119764 260176 119770 260188
rect 144914 260176 144920 260188
rect 144972 260176 144978 260228
rect 145006 260176 145012 260228
rect 145064 260216 145070 260228
rect 146248 260216 146254 260228
rect 145064 260188 146254 260216
rect 145064 260176 145070 260188
rect 146248 260176 146254 260188
rect 146306 260176 146312 260228
rect 147674 260176 147680 260228
rect 147732 260216 147738 260228
rect 148732 260216 148738 260228
rect 147732 260188 148738 260216
rect 147732 260176 147738 260188
rect 148732 260176 148738 260188
rect 148790 260176 148796 260228
rect 149054 260176 149060 260228
rect 149112 260216 149118 260228
rect 190546 260216 190552 260228
rect 149112 260188 190552 260216
rect 149112 260176 149118 260188
rect 190546 260176 190552 260188
rect 190604 260176 190610 260228
rect 115474 260108 115480 260160
rect 115532 260148 115538 260160
rect 129734 260148 129740 260160
rect 115532 260120 129740 260148
rect 115532 260108 115538 260120
rect 129734 260108 129740 260120
rect 129792 260108 129798 260160
rect 142154 260108 142160 260160
rect 142212 260148 142218 260160
rect 192294 260148 192300 260160
rect 142212 260120 192300 260148
rect 142212 260108 142218 260120
rect 192294 260108 192300 260120
rect 192352 260108 192358 260160
rect 120166 260040 120172 260092
rect 120224 260080 120230 260092
rect 121362 260080 121368 260092
rect 120224 260052 121368 260080
rect 120224 260040 120230 260052
rect 121362 260040 121368 260052
rect 121420 260040 121426 260092
rect 160094 260040 160100 260092
rect 160152 260080 160158 260092
rect 161152 260080 161158 260092
rect 160152 260052 161158 260080
rect 160152 260040 160158 260052
rect 161152 260040 161158 260052
rect 161210 260040 161216 260092
rect 178034 260040 178040 260092
rect 178092 260080 178098 260092
rect 179368 260080 179374 260092
rect 178092 260052 179374 260080
rect 178092 260040 178098 260052
rect 179368 260040 179374 260052
rect 179426 260040 179432 260092
rect 192018 260080 192024 260092
rect 180766 260052 192024 260080
rect 115198 259972 115204 260024
rect 115256 260012 115262 260024
rect 126054 260012 126060 260024
rect 115256 259984 126060 260012
rect 115256 259972 115262 259984
rect 126054 259972 126060 259984
rect 126112 259972 126118 260024
rect 180334 259972 180340 260024
rect 180392 260012 180398 260024
rect 180766 260012 180794 260052
rect 192018 260040 192024 260052
rect 192076 260040 192082 260092
rect 180392 259984 180794 260012
rect 180392 259972 180398 259984
rect 184658 259972 184664 260024
rect 184716 260012 184722 260024
rect 196434 260012 196440 260024
rect 184716 259984 196440 260012
rect 184716 259972 184722 259984
rect 196434 259972 196440 259984
rect 196492 259972 196498 260024
rect 114002 259904 114008 259956
rect 114060 259944 114066 259956
rect 123202 259944 123208 259956
rect 114060 259916 123208 259944
rect 114060 259904 114066 259916
rect 123202 259904 123208 259916
rect 123260 259944 123266 259956
rect 123570 259944 123576 259956
rect 123260 259916 123576 259944
rect 123260 259904 123266 259916
rect 123570 259904 123576 259916
rect 123628 259904 123634 259956
rect 178862 259904 178868 259956
rect 178920 259944 178926 259956
rect 197722 259944 197728 259956
rect 178920 259916 197728 259944
rect 178920 259904 178926 259916
rect 197722 259904 197728 259916
rect 197780 259904 197786 259956
rect 116670 259836 116676 259888
rect 116728 259876 116734 259888
rect 128446 259876 128452 259888
rect 116728 259848 128452 259876
rect 116728 259836 116734 259848
rect 128446 259836 128452 259848
rect 128504 259836 128510 259888
rect 179506 259836 179512 259888
rect 179564 259876 179570 259888
rect 197906 259876 197912 259888
rect 179564 259848 197912 259876
rect 179564 259836 179570 259848
rect 197906 259836 197912 259848
rect 197964 259836 197970 259888
rect 112530 259768 112536 259820
rect 112588 259808 112594 259820
rect 131114 259808 131120 259820
rect 112588 259780 131120 259808
rect 112588 259768 112594 259780
rect 131114 259768 131120 259780
rect 131172 259768 131178 259820
rect 167914 259768 167920 259820
rect 167972 259808 167978 259820
rect 192202 259808 192208 259820
rect 167972 259780 192208 259808
rect 167972 259768 167978 259780
rect 192202 259768 192208 259780
rect 192260 259768 192266 259820
rect 115382 259700 115388 259752
rect 115440 259740 115446 259752
rect 145006 259740 145012 259752
rect 115440 259712 145012 259740
rect 115440 259700 115446 259712
rect 145006 259700 145012 259712
rect 145064 259700 145070 259752
rect 172238 259700 172244 259752
rect 172296 259740 172302 259752
rect 197814 259740 197820 259752
rect 172296 259712 197820 259740
rect 172296 259700 172302 259712
rect 197814 259700 197820 259712
rect 197872 259700 197878 259752
rect 116762 259632 116768 259684
rect 116820 259672 116826 259684
rect 147674 259672 147680 259684
rect 116820 259644 147680 259672
rect 116820 259632 116826 259644
rect 147674 259632 147680 259644
rect 147732 259632 147738 259684
rect 166442 259632 166448 259684
rect 166500 259672 166506 259684
rect 197078 259672 197084 259684
rect 166500 259644 197084 259672
rect 166500 259632 166506 259644
rect 197078 259632 197084 259644
rect 197136 259632 197142 259684
rect 113910 259564 113916 259616
rect 113968 259604 113974 259616
rect 146754 259604 146760 259616
rect 113968 259576 146760 259604
rect 113968 259564 113974 259576
rect 146754 259564 146760 259576
rect 146812 259564 146818 259616
rect 162302 259564 162308 259616
rect 162360 259604 162366 259616
rect 195238 259604 195244 259616
rect 162360 259576 195244 259604
rect 162360 259564 162366 259576
rect 195238 259564 195244 259576
rect 195296 259564 195302 259616
rect 116578 259496 116584 259548
rect 116636 259536 116642 259548
rect 149146 259536 149152 259548
rect 116636 259508 149152 259536
rect 116636 259496 116642 259508
rect 149146 259496 149152 259508
rect 149204 259496 149210 259548
rect 175366 259496 175372 259548
rect 175424 259536 175430 259548
rect 192110 259536 192116 259548
rect 175424 259508 192116 259536
rect 175424 259496 175430 259508
rect 192110 259496 192116 259508
rect 192168 259496 192174 259548
rect 117866 259428 117872 259480
rect 117924 259468 117930 259480
rect 150894 259468 150900 259480
rect 117924 259440 150900 259468
rect 117924 259428 117930 259440
rect 150894 259428 150900 259440
rect 150952 259428 150958 259480
rect 176378 259428 176384 259480
rect 176436 259468 176442 259480
rect 195054 259468 195060 259480
rect 176436 259440 195060 259468
rect 176436 259428 176442 259440
rect 195054 259428 195060 259440
rect 195112 259428 195118 259480
rect 3234 256708 3240 256760
rect 3292 256748 3298 256760
rect 117314 256748 117320 256760
rect 3292 256720 117320 256748
rect 3292 256708 3298 256720
rect 117314 256708 117320 256720
rect 117372 256708 117378 256760
rect 191650 253920 191656 253972
rect 191708 253960 191714 253972
rect 579798 253960 579804 253972
rect 191708 253932 579804 253960
rect 191708 253920 191714 253932
rect 579798 253920 579804 253932
rect 579856 253920 579862 253972
rect 120074 253172 120080 253224
rect 120132 253212 120138 253224
rect 120350 253212 120356 253224
rect 120132 253184 120356 253212
rect 120132 253172 120138 253184
rect 120350 253172 120356 253184
rect 120408 253172 120414 253224
rect 3142 252560 3148 252612
rect 3200 252600 3206 252612
rect 119338 252600 119344 252612
rect 3200 252572 119344 252600
rect 3200 252560 3206 252572
rect 119338 252560 119344 252572
rect 119396 252560 119402 252612
rect 192570 251132 192576 251184
rect 192628 251172 192634 251184
rect 579982 251172 579988 251184
rect 192628 251144 579988 251172
rect 192628 251132 192634 251144
rect 579982 251132 579988 251144
rect 580040 251132 580046 251184
rect 191190 241476 191196 241528
rect 191248 241516 191254 241528
rect 580166 241516 580172 241528
rect 191248 241488 580172 241516
rect 191248 241476 191254 241488
rect 580166 241476 580172 241488
rect 580224 241476 580230 241528
rect 3326 240116 3332 240168
rect 3384 240156 3390 240168
rect 119430 240156 119436 240168
rect 3384 240128 119436 240156
rect 3384 240116 3390 240128
rect 119430 240116 119436 240128
rect 119488 240116 119494 240168
rect 498838 238688 498844 238740
rect 498896 238728 498902 238740
rect 580166 238728 580172 238740
rect 498896 238700 580172 238728
rect 498896 238688 498902 238700
rect 580166 238688 580172 238700
rect 580224 238688 580230 238740
rect 3326 229100 3332 229152
rect 3384 229140 3390 229152
rect 120902 229140 120908 229152
rect 3384 229112 120908 229140
rect 3384 229100 3390 229112
rect 120902 229100 120908 229112
rect 120960 229100 120966 229152
rect 190086 224952 190092 225004
rect 190144 224992 190150 225004
rect 579982 224992 579988 225004
rect 190144 224964 579988 224992
rect 190144 224952 190150 224964
rect 579982 224952 579988 224964
rect 580040 224952 580046 225004
rect 3050 220804 3056 220856
rect 3108 220844 3114 220856
rect 119522 220844 119528 220856
rect 3108 220816 119528 220844
rect 3108 220804 3114 220816
rect 119522 220804 119528 220816
rect 119580 220804 119586 220856
rect 3142 208360 3148 208412
rect 3200 208400 3206 208412
rect 120534 208400 120540 208412
rect 3200 208372 120540 208400
rect 3200 208360 3206 208372
rect 120534 208360 120540 208372
rect 120592 208360 120598 208412
rect 190546 204892 190552 204944
rect 190604 204932 190610 204944
rect 190914 204932 190920 204944
rect 190604 204904 190920 204932
rect 190604 204892 190610 204904
rect 190914 204892 190920 204904
rect 190972 204892 190978 204944
rect 96062 201492 96068 201544
rect 96120 201532 96126 201544
rect 118694 201532 118700 201544
rect 96120 201504 118700 201532
rect 96120 201492 96126 201504
rect 118694 201492 118700 201504
rect 118752 201532 118758 201544
rect 118970 201532 118976 201544
rect 118752 201504 118976 201532
rect 118752 201492 118758 201504
rect 118970 201492 118976 201504
rect 119028 201492 119034 201544
rect 191466 201492 191472 201544
rect 191524 201532 191530 201544
rect 191742 201532 191748 201544
rect 191524 201504 191748 201532
rect 191524 201492 191530 201504
rect 191742 201492 191748 201504
rect 191800 201532 191806 201544
rect 204254 201532 204260 201544
rect 191800 201504 204260 201532
rect 191800 201492 191806 201504
rect 204254 201492 204260 201504
rect 204312 201492 204318 201544
rect 115934 201424 115940 201476
rect 115992 201464 115998 201476
rect 117038 201464 117044 201476
rect 115992 201436 117044 201464
rect 115992 201424 115998 201436
rect 117038 201424 117044 201436
rect 117096 201424 117102 201476
rect 3602 200812 3608 200864
rect 3660 200852 3666 200864
rect 95142 200852 95148 200864
rect 3660 200824 95148 200852
rect 3660 200812 3666 200824
rect 95142 200812 95148 200824
rect 95200 200812 95206 200864
rect 96246 200812 96252 200864
rect 96304 200852 96310 200864
rect 117314 200852 117320 200864
rect 96304 200824 117320 200852
rect 96304 200812 96310 200824
rect 117314 200812 117320 200824
rect 117372 200852 117378 200864
rect 117372 200824 121040 200852
rect 117372 200812 117378 200824
rect 3510 200744 3516 200796
rect 3568 200784 3574 200796
rect 96430 200784 96436 200796
rect 3568 200756 96436 200784
rect 3568 200744 3574 200756
rect 96430 200744 96436 200756
rect 96488 200744 96494 200796
rect 109954 200744 109960 200796
rect 110012 200784 110018 200796
rect 110012 200756 118004 200784
rect 110012 200744 110018 200756
rect 104526 200472 104532 200524
rect 104584 200512 104590 200524
rect 113174 200512 113180 200524
rect 104584 200484 113180 200512
rect 104584 200472 104590 200484
rect 113174 200472 113180 200484
rect 113232 200472 113238 200524
rect 117976 200512 118004 200756
rect 121012 200716 121040 200824
rect 204346 200812 204352 200864
rect 204404 200852 204410 200864
rect 252554 200852 252560 200864
rect 204404 200824 252560 200852
rect 204404 200812 204410 200824
rect 252554 200812 252560 200824
rect 252612 200812 252618 200864
rect 121178 200744 121184 200796
rect 121236 200784 121242 200796
rect 580718 200784 580724 200796
rect 121236 200756 125732 200784
rect 121236 200744 121242 200756
rect 125704 200728 125732 200756
rect 128326 200756 167868 200784
rect 125548 200716 125554 200728
rect 121012 200688 125554 200716
rect 125548 200676 125554 200688
rect 125606 200676 125612 200728
rect 125686 200676 125692 200728
rect 125744 200676 125750 200728
rect 119522 200608 119528 200660
rect 119580 200648 119586 200660
rect 128326 200648 128354 200756
rect 142126 200688 143534 200716
rect 142126 200648 142154 200688
rect 119580 200620 128354 200648
rect 129706 200620 142154 200648
rect 143506 200648 143534 200688
rect 144886 200688 161566 200716
rect 144886 200648 144914 200688
rect 143506 200620 144914 200648
rect 119580 200608 119586 200620
rect 119338 200540 119344 200592
rect 119396 200580 119402 200592
rect 129706 200580 129734 200620
rect 119396 200552 129734 200580
rect 119396 200540 119402 200552
rect 132126 200540 132132 200592
rect 132184 200580 132190 200592
rect 132184 200552 141970 200580
rect 132184 200540 132190 200552
rect 121178 200512 121184 200524
rect 117976 200484 121184 200512
rect 121178 200472 121184 200484
rect 121236 200472 121242 200524
rect 124398 200472 124404 200524
rect 124456 200512 124462 200524
rect 131758 200512 131764 200524
rect 124456 200484 131764 200512
rect 124456 200472 124462 200484
rect 131758 200472 131764 200484
rect 131816 200472 131822 200524
rect 131850 200472 131856 200524
rect 131908 200512 131914 200524
rect 131908 200484 141878 200512
rect 131908 200472 131914 200484
rect 104434 200404 104440 200456
rect 104492 200444 104498 200456
rect 118786 200444 118792 200456
rect 104492 200416 118792 200444
rect 104492 200404 104498 200416
rect 118786 200404 118792 200416
rect 118844 200404 118850 200456
rect 120534 200404 120540 200456
rect 120592 200444 120598 200456
rect 120994 200444 121000 200456
rect 120592 200416 121000 200444
rect 120592 200404 120598 200416
rect 120994 200404 121000 200416
rect 121052 200404 121058 200456
rect 124186 200416 135254 200444
rect 97534 200336 97540 200388
rect 97592 200376 97598 200388
rect 115934 200376 115940 200388
rect 97592 200348 115940 200376
rect 97592 200336 97598 200348
rect 115934 200336 115940 200348
rect 115992 200336 115998 200388
rect 94958 200268 94964 200320
rect 95016 200308 95022 200320
rect 120258 200308 120264 200320
rect 95016 200280 120264 200308
rect 95016 200268 95022 200280
rect 120258 200268 120264 200280
rect 120316 200268 120322 200320
rect 123202 200268 123208 200320
rect 123260 200308 123266 200320
rect 124186 200308 124214 200416
rect 132126 200308 132132 200320
rect 123260 200280 124214 200308
rect 128326 200280 132132 200308
rect 123260 200268 123266 200280
rect 96430 200200 96436 200252
rect 96488 200240 96494 200252
rect 128326 200240 128354 200280
rect 132126 200268 132132 200280
rect 132184 200268 132190 200320
rect 135226 200308 135254 200416
rect 135226 200280 137922 200308
rect 96488 200212 128354 200240
rect 96488 200200 96494 200212
rect 132034 200200 132040 200252
rect 132092 200240 132098 200252
rect 132092 200212 135254 200240
rect 132092 200200 132098 200212
rect 95142 200132 95148 200184
rect 95200 200172 95206 200184
rect 131850 200172 131856 200184
rect 95200 200144 131856 200172
rect 95200 200132 95206 200144
rect 131850 200132 131856 200144
rect 131908 200132 131914 200184
rect 131942 200132 131948 200184
rect 132000 200172 132006 200184
rect 135226 200172 135254 200212
rect 132000 200144 133874 200172
rect 135226 200144 135990 200172
rect 132000 200132 132006 200144
rect 133846 200104 133874 200144
rect 135962 200104 135990 200144
rect 133846 200076 135898 200104
rect 135962 200076 136174 200104
rect 129734 199996 129740 200048
rect 129792 200036 129798 200048
rect 129792 200008 134058 200036
rect 129792 199996 129798 200008
rect 131850 199928 131856 199980
rect 131908 199968 131914 199980
rect 131908 199940 132770 199968
rect 131908 199928 131914 199940
rect 132218 199900 132224 199912
rect 124186 199872 132224 199900
rect 120994 199792 121000 199844
rect 121052 199832 121058 199844
rect 124186 199832 124214 199872
rect 132218 199860 132224 199872
rect 132276 199860 132282 199912
rect 132632 199860 132638 199912
rect 132690 199860 132696 199912
rect 121052 199804 124214 199832
rect 121052 199792 121058 199804
rect 127894 199792 127900 199844
rect 127952 199832 127958 199844
rect 127952 199804 130516 199832
rect 127952 199792 127958 199804
rect 119338 199724 119344 199776
rect 119396 199764 119402 199776
rect 130488 199764 130516 199804
rect 131850 199792 131856 199844
rect 131908 199832 131914 199844
rect 132650 199832 132678 199860
rect 132742 199844 132770 199940
rect 134030 199912 134058 200008
rect 133000 199860 133006 199912
rect 133058 199860 133064 199912
rect 133092 199860 133098 199912
rect 133150 199860 133156 199912
rect 133800 199872 133966 199900
rect 131908 199804 132678 199832
rect 131908 199792 131914 199804
rect 132724 199792 132730 199844
rect 132782 199792 132788 199844
rect 133018 199764 133046 199860
rect 119396 199736 130424 199764
rect 130488 199736 133046 199764
rect 133110 199776 133138 199860
rect 133110 199736 133144 199776
rect 119396 199724 119402 199736
rect 84194 199520 84200 199572
rect 84252 199560 84258 199572
rect 128446 199560 128452 199572
rect 84252 199532 128452 199560
rect 84252 199520 84258 199532
rect 128446 199520 128452 199532
rect 128504 199560 128510 199572
rect 129642 199560 129648 199572
rect 128504 199532 129648 199560
rect 128504 199520 128510 199532
rect 129642 199520 129648 199532
rect 129700 199520 129706 199572
rect 130396 199560 130424 199736
rect 133138 199724 133144 199736
rect 133196 199724 133202 199776
rect 133800 199764 133828 199872
rect 133248 199736 133828 199764
rect 131758 199656 131764 199708
rect 131816 199696 131822 199708
rect 133248 199696 133276 199736
rect 133782 199696 133788 199708
rect 131816 199668 133276 199696
rect 133708 199668 133788 199696
rect 131816 199656 131822 199668
rect 133708 199640 133736 199668
rect 133782 199656 133788 199668
rect 133840 199656 133846 199708
rect 133938 199696 133966 199872
rect 134012 199860 134018 199912
rect 134070 199860 134076 199912
rect 134104 199860 134110 199912
rect 134162 199860 134168 199912
rect 134564 199900 134570 199912
rect 134536 199860 134570 199900
rect 134622 199860 134628 199912
rect 134932 199860 134938 199912
rect 134990 199860 134996 199912
rect 135392 199900 135398 199912
rect 135272 199872 135398 199900
rect 134122 199776 134150 199860
rect 134122 199736 134156 199776
rect 134150 199724 134156 199736
rect 134208 199724 134214 199776
rect 134058 199696 134064 199708
rect 133938 199668 134064 199696
rect 134058 199656 134064 199668
rect 134116 199656 134122 199708
rect 134536 199640 134564 199860
rect 134950 199640 134978 199860
rect 133690 199588 133696 199640
rect 133748 199588 133754 199640
rect 134518 199588 134524 199640
rect 134576 199588 134582 199640
rect 134886 199588 134892 199640
rect 134944 199600 134978 199640
rect 134944 199588 134950 199600
rect 131666 199560 131672 199572
rect 130396 199532 131672 199560
rect 131666 199520 131672 199532
rect 131724 199520 131730 199572
rect 131850 199520 131856 199572
rect 131908 199560 131914 199572
rect 133598 199560 133604 199572
rect 131908 199532 133604 199560
rect 131908 199520 131914 199532
rect 133598 199520 133604 199532
rect 133656 199520 133662 199572
rect 133782 199520 133788 199572
rect 133840 199560 133846 199572
rect 134334 199560 134340 199572
rect 133840 199532 134340 199560
rect 133840 199520 133846 199532
rect 134334 199520 134340 199532
rect 134392 199520 134398 199572
rect 135272 199560 135300 199872
rect 135392 199860 135398 199872
rect 135450 199860 135456 199912
rect 135760 199860 135766 199912
rect 135818 199860 135824 199912
rect 135778 199832 135806 199860
rect 135364 199804 135806 199832
rect 135364 199628 135392 199804
rect 135714 199628 135720 199640
rect 135364 199600 135720 199628
rect 135714 199588 135720 199600
rect 135772 199588 135778 199640
rect 135346 199560 135352 199572
rect 135272 199532 135352 199560
rect 135346 199520 135352 199532
rect 135404 199520 135410 199572
rect 135870 199560 135898 200076
rect 136146 199912 136174 200076
rect 136836 199940 137738 199968
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136128 199860 136134 199912
rect 136186 199860 136192 199912
rect 136220 199860 136226 199912
rect 136278 199860 136284 199912
rect 136404 199860 136410 199912
rect 136462 199860 136468 199912
rect 136836 199900 136864 199940
rect 137710 199912 137738 199940
rect 136560 199872 136864 199900
rect 136054 199776 136082 199860
rect 136238 199776 136266 199860
rect 136054 199736 136088 199776
rect 136082 199724 136088 199736
rect 136140 199724 136146 199776
rect 136174 199724 136180 199776
rect 136232 199736 136266 199776
rect 136232 199724 136238 199736
rect 136422 199708 136450 199860
rect 136422 199668 136456 199708
rect 136450 199656 136456 199668
rect 136508 199656 136514 199708
rect 136358 199588 136364 199640
rect 136416 199628 136422 199640
rect 136560 199628 136588 199872
rect 137232 199860 137238 199912
rect 137290 199900 137296 199912
rect 137290 199872 137508 199900
rect 137290 199860 137296 199872
rect 136680 199792 136686 199844
rect 136738 199792 136744 199844
rect 137140 199792 137146 199844
rect 137198 199832 137204 199844
rect 137198 199792 137232 199832
rect 137324 199792 137330 199844
rect 137382 199792 137388 199844
rect 136416 199600 136588 199628
rect 136416 199588 136422 199600
rect 136698 199560 136726 199792
rect 137204 199708 137232 199792
rect 137342 199708 137370 199792
rect 137186 199656 137192 199708
rect 137244 199656 137250 199708
rect 137278 199656 137284 199708
rect 137336 199668 137370 199708
rect 137336 199656 137342 199668
rect 137480 199572 137508 199872
rect 137600 199860 137606 199912
rect 137658 199860 137664 199912
rect 137692 199860 137698 199912
rect 137750 199860 137756 199912
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 137618 199776 137646 199860
rect 137618 199736 137652 199776
rect 137646 199724 137652 199736
rect 137704 199724 137710 199776
rect 137802 199708 137830 199860
rect 137738 199656 137744 199708
rect 137796 199668 137830 199708
rect 137796 199656 137802 199668
rect 137894 199640 137922 200280
rect 139550 199940 140498 199968
rect 137968 199860 137974 199912
rect 138026 199860 138032 199912
rect 138704 199860 138710 199912
rect 138762 199860 138768 199912
rect 138796 199860 138802 199912
rect 138854 199860 138860 199912
rect 138888 199860 138894 199912
rect 138946 199860 138952 199912
rect 139164 199860 139170 199912
rect 139222 199860 139228 199912
rect 139440 199900 139446 199912
rect 139412 199860 139446 199900
rect 139498 199860 139504 199912
rect 137830 199588 137836 199640
rect 137888 199600 137922 199640
rect 137888 199588 137894 199600
rect 135870 199532 136726 199560
rect 137462 199520 137468 199572
rect 137520 199520 137526 199572
rect 137986 199560 138014 199860
rect 138290 199560 138296 199572
rect 137986 199532 138296 199560
rect 138290 199520 138296 199532
rect 138348 199520 138354 199572
rect 138474 199520 138480 199572
rect 138532 199560 138538 199572
rect 138722 199560 138750 199860
rect 138814 199776 138842 199860
rect 138906 199832 138934 199860
rect 138906 199804 138980 199832
rect 138814 199736 138848 199776
rect 138842 199724 138848 199736
rect 138900 199724 138906 199776
rect 138532 199532 138750 199560
rect 138532 199520 138538 199532
rect 138842 199520 138848 199572
rect 138900 199560 138906 199572
rect 138952 199560 138980 199804
rect 139182 199640 139210 199860
rect 139412 199776 139440 199860
rect 139394 199724 139400 199776
rect 139452 199724 139458 199776
rect 139550 199640 139578 199940
rect 140470 199912 140498 199940
rect 140562 199940 141234 199968
rect 139716 199860 139722 199912
rect 139774 199860 139780 199912
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 140452 199860 140458 199912
rect 140510 199860 140516 199912
rect 139734 199640 139762 199860
rect 139918 199696 139946 199860
rect 140562 199832 140590 199940
rect 141206 199912 141234 199940
rect 140636 199860 140642 199912
rect 140694 199860 140700 199912
rect 140820 199860 140826 199912
rect 140878 199860 140884 199912
rect 141096 199860 141102 199912
rect 141154 199860 141160 199912
rect 141188 199860 141194 199912
rect 141246 199860 141252 199912
rect 141280 199860 141286 199912
rect 141338 199860 141344 199912
rect 141372 199860 141378 199912
rect 141430 199900 141436 199912
rect 141430 199860 141464 199900
rect 139872 199668 139946 199696
rect 140332 199804 140590 199832
rect 139872 199640 139900 199668
rect 140332 199640 140360 199804
rect 140654 199696 140682 199860
rect 140838 199764 140866 199860
rect 140838 199736 141004 199764
rect 140516 199668 140682 199696
rect 139118 199588 139124 199640
rect 139176 199600 139210 199640
rect 139176 199588 139182 199600
rect 139486 199588 139492 199640
rect 139544 199600 139578 199640
rect 139544 199588 139550 199600
rect 139670 199588 139676 199640
rect 139728 199600 139762 199640
rect 139728 199588 139734 199600
rect 139854 199588 139860 199640
rect 139912 199588 139918 199640
rect 140314 199588 140320 199640
rect 140372 199588 140378 199640
rect 138900 199532 138980 199560
rect 140056 199532 140360 199560
rect 138900 199520 138906 199532
rect 46934 199452 46940 199504
rect 46992 199492 46998 199504
rect 138934 199492 138940 199504
rect 46992 199464 138940 199492
rect 46992 199452 46998 199464
rect 138934 199452 138940 199464
rect 138992 199452 138998 199504
rect 4062 199384 4068 199436
rect 4120 199424 4126 199436
rect 140056 199424 140084 199532
rect 4120 199396 140084 199424
rect 4120 199384 4126 199396
rect 121270 199316 121276 199368
rect 121328 199356 121334 199368
rect 140038 199356 140044 199368
rect 121328 199328 140044 199356
rect 121328 199316 121334 199328
rect 140038 199316 140044 199328
rect 140096 199316 140102 199368
rect 140332 199356 140360 199532
rect 140516 199424 140544 199668
rect 140976 199640 141004 199736
rect 141114 199708 141142 199860
rect 141298 199776 141326 199860
rect 141234 199724 141240 199776
rect 141292 199736 141326 199776
rect 141292 199724 141298 199736
rect 141114 199668 141148 199708
rect 141142 199656 141148 199668
rect 141200 199656 141206 199708
rect 141326 199656 141332 199708
rect 141384 199696 141390 199708
rect 141436 199696 141464 199860
rect 141384 199668 141464 199696
rect 141384 199656 141390 199668
rect 140958 199588 140964 199640
rect 141016 199588 141022 199640
rect 141050 199588 141056 199640
rect 141108 199628 141114 199640
rect 141510 199628 141516 199640
rect 141108 199600 141516 199628
rect 141108 199588 141114 199600
rect 141510 199588 141516 199600
rect 141568 199588 141574 199640
rect 141850 199560 141878 200484
rect 141942 199912 141970 200552
rect 159284 200552 160094 200580
rect 144886 200484 150802 200512
rect 144886 200308 144914 200484
rect 143092 200280 144914 200308
rect 144978 200416 149744 200444
rect 141924 199860 141930 199912
rect 141982 199860 141988 199912
rect 142200 199860 142206 199912
rect 142258 199860 142264 199912
rect 142292 199860 142298 199912
rect 142350 199860 142356 199912
rect 142384 199860 142390 199912
rect 142442 199900 142448 199912
rect 142442 199860 142476 199900
rect 142568 199860 142574 199912
rect 142626 199860 142632 199912
rect 142660 199860 142666 199912
rect 142718 199860 142724 199912
rect 142752 199860 142758 199912
rect 142810 199860 142816 199912
rect 142844 199860 142850 199912
rect 142902 199860 142908 199912
rect 142218 199776 142246 199860
rect 142154 199724 142160 199776
rect 142212 199736 142246 199776
rect 142212 199724 142218 199736
rect 142310 199708 142338 199860
rect 142448 199776 142476 199860
rect 142586 199832 142614 199860
rect 142540 199804 142614 199832
rect 142430 199724 142436 199776
rect 142488 199724 142494 199776
rect 142540 199708 142568 199804
rect 142678 199776 142706 199860
rect 142614 199724 142620 199776
rect 142672 199736 142706 199776
rect 142672 199724 142678 199736
rect 142770 199708 142798 199860
rect 142862 199776 142890 199860
rect 142862 199736 142896 199776
rect 142890 199724 142896 199736
rect 142948 199724 142954 199776
rect 142246 199656 142252 199708
rect 142304 199668 142338 199708
rect 142304 199656 142310 199668
rect 142522 199656 142528 199708
rect 142580 199656 142586 199708
rect 142706 199656 142712 199708
rect 142764 199668 142798 199708
rect 142764 199656 142770 199668
rect 143092 199640 143120 200280
rect 144978 200240 145006 200416
rect 144886 200212 145006 200240
rect 144886 200036 144914 200212
rect 144150 200008 144914 200036
rect 147646 200076 148410 200104
rect 143488 199860 143494 199912
rect 143546 199860 143552 199912
rect 143764 199860 143770 199912
rect 143822 199860 143828 199912
rect 144040 199860 144046 199912
rect 144098 199860 144104 199912
rect 143074 199588 143080 199640
rect 143132 199588 143138 199640
rect 142430 199560 142436 199572
rect 141850 199532 142436 199560
rect 142430 199520 142436 199532
rect 142488 199520 142494 199572
rect 143506 199504 143534 199860
rect 143782 199572 143810 199860
rect 144058 199572 144086 199860
rect 143718 199520 143724 199572
rect 143776 199532 143810 199572
rect 143776 199520 143782 199532
rect 143994 199520 144000 199572
rect 144052 199532 144086 199572
rect 144052 199520 144058 199532
rect 144150 199504 144178 200008
rect 147646 199968 147674 200076
rect 144564 199940 146064 199968
rect 144316 199860 144322 199912
rect 144374 199860 144380 199912
rect 144334 199696 144362 199860
rect 144334 199668 144500 199696
rect 144472 199640 144500 199668
rect 144454 199588 144460 199640
rect 144512 199588 144518 199640
rect 141050 199452 141056 199504
rect 141108 199492 141114 199504
rect 142706 199492 142712 199504
rect 141108 199464 142712 199492
rect 141108 199452 141114 199464
rect 142706 199452 142712 199464
rect 142764 199452 142770 199504
rect 143442 199452 143448 199504
rect 143500 199464 143534 199504
rect 143500 199452 143506 199464
rect 144086 199452 144092 199504
rect 144144 199464 144178 199504
rect 144144 199452 144150 199464
rect 140590 199424 140596 199436
rect 140516 199396 140596 199424
rect 140590 199384 140596 199396
rect 140648 199384 140654 199436
rect 140774 199384 140780 199436
rect 140832 199424 140838 199436
rect 144564 199424 144592 199940
rect 144684 199860 144690 199912
rect 144742 199860 144748 199912
rect 144776 199860 144782 199912
rect 144834 199860 144840 199912
rect 145052 199860 145058 199912
rect 145110 199860 145116 199912
rect 145420 199900 145426 199912
rect 145392 199860 145426 199900
rect 145478 199860 145484 199912
rect 145512 199860 145518 199912
rect 145570 199860 145576 199912
rect 145604 199860 145610 199912
rect 145662 199860 145668 199912
rect 145880 199860 145886 199912
rect 145938 199860 145944 199912
rect 144702 199764 144730 199860
rect 144656 199736 144730 199764
rect 144656 199572 144684 199736
rect 144794 199708 144822 199860
rect 144730 199656 144736 199708
rect 144788 199668 144822 199708
rect 144788 199656 144794 199668
rect 145070 199572 145098 199860
rect 145236 199792 145242 199844
rect 145294 199792 145300 199844
rect 144638 199520 144644 199572
rect 144696 199520 144702 199572
rect 145006 199520 145012 199572
rect 145064 199532 145098 199572
rect 145064 199520 145070 199532
rect 144730 199452 144736 199504
rect 144788 199492 144794 199504
rect 145254 199492 145282 199792
rect 145392 199640 145420 199860
rect 145530 199832 145558 199860
rect 145484 199804 145558 199832
rect 145484 199708 145512 199804
rect 145622 199708 145650 199860
rect 145466 199656 145472 199708
rect 145524 199656 145530 199708
rect 145558 199656 145564 199708
rect 145616 199668 145650 199708
rect 145616 199656 145622 199668
rect 145374 199588 145380 199640
rect 145432 199588 145438 199640
rect 144788 199464 145282 199492
rect 144788 199452 144794 199464
rect 140832 199396 144592 199424
rect 140832 199384 140838 199396
rect 145898 199368 145926 199860
rect 146036 199492 146064 199940
rect 147508 199940 147674 199968
rect 147830 200008 148318 200036
rect 146248 199860 146254 199912
rect 146306 199860 146312 199912
rect 146340 199860 146346 199912
rect 146398 199860 146404 199912
rect 146524 199860 146530 199912
rect 146582 199860 146588 199912
rect 146800 199860 146806 199912
rect 146858 199860 146864 199912
rect 146892 199860 146898 199912
rect 146950 199860 146956 199912
rect 147168 199900 147174 199912
rect 147140 199860 147174 199900
rect 147226 199860 147232 199912
rect 147260 199860 147266 199912
rect 147318 199860 147324 199912
rect 146266 199572 146294 199860
rect 146358 199640 146386 199860
rect 146542 199708 146570 199860
rect 146616 199792 146622 199844
rect 146674 199792 146680 199844
rect 146478 199656 146484 199708
rect 146536 199668 146570 199708
rect 146634 199708 146662 199792
rect 146634 199668 146668 199708
rect 146536 199656 146542 199668
rect 146662 199656 146668 199668
rect 146720 199656 146726 199708
rect 146818 199640 146846 199860
rect 146910 199708 146938 199860
rect 146984 199792 146990 199844
rect 147042 199832 147048 199844
rect 147042 199792 147076 199832
rect 146910 199668 146944 199708
rect 146938 199656 146944 199668
rect 146996 199656 147002 199708
rect 146358 199600 146392 199640
rect 146386 199588 146392 199600
rect 146444 199588 146450 199640
rect 146754 199588 146760 199640
rect 146812 199600 146846 199640
rect 146812 199588 146818 199600
rect 146266 199532 146300 199572
rect 146294 199520 146300 199532
rect 146352 199520 146358 199572
rect 146570 199520 146576 199572
rect 146628 199560 146634 199572
rect 147048 199560 147076 199792
rect 146628 199532 147076 199560
rect 146628 199520 146634 199532
rect 146036 199464 146294 199492
rect 146266 199424 146294 199464
rect 147140 199424 147168 199860
rect 147278 199640 147306 199860
rect 147508 199640 147536 199940
rect 147628 199900 147634 199912
rect 147600 199860 147634 199900
rect 147686 199860 147692 199912
rect 147720 199860 147726 199912
rect 147778 199860 147784 199912
rect 147214 199588 147220 199640
rect 147272 199600 147306 199640
rect 147272 199588 147278 199600
rect 147490 199588 147496 199640
rect 147548 199588 147554 199640
rect 146266 199396 147168 199424
rect 140332 199328 145788 199356
rect 107562 199248 107568 199300
rect 107620 199288 107626 199300
rect 133598 199288 133604 199300
rect 107620 199260 133604 199288
rect 107620 199248 107626 199260
rect 133598 199248 133604 199260
rect 133656 199248 133662 199300
rect 135070 199248 135076 199300
rect 135128 199288 135134 199300
rect 135622 199288 135628 199300
rect 135128 199260 135628 199288
rect 135128 199248 135134 199260
rect 135622 199248 135628 199260
rect 135680 199248 135686 199300
rect 138014 199248 138020 199300
rect 138072 199288 138078 199300
rect 145650 199288 145656 199300
rect 138072 199260 145656 199288
rect 138072 199248 138078 199260
rect 145650 199248 145656 199260
rect 145708 199248 145714 199300
rect 129642 199180 129648 199232
rect 129700 199220 129706 199232
rect 141418 199220 141424 199232
rect 129700 199192 141424 199220
rect 129700 199180 129706 199192
rect 141418 199180 141424 199192
rect 141476 199180 141482 199232
rect 145760 199220 145788 199328
rect 145834 199316 145840 199368
rect 145892 199328 145926 199368
rect 145892 199316 145898 199328
rect 146570 199248 146576 199300
rect 146628 199288 146634 199300
rect 147600 199288 147628 199860
rect 147738 199708 147766 199860
rect 147674 199656 147680 199708
rect 147732 199668 147766 199708
rect 147732 199656 147738 199668
rect 147830 199640 147858 200008
rect 147922 199940 148226 199968
rect 147922 199912 147950 199940
rect 147904 199860 147910 199912
rect 147962 199860 147968 199912
rect 147996 199860 148002 199912
rect 148054 199860 148060 199912
rect 148088 199860 148094 199912
rect 148146 199860 148152 199912
rect 148014 199776 148042 199860
rect 147950 199724 147956 199776
rect 148008 199736 148042 199776
rect 148008 199724 148014 199736
rect 148106 199696 148134 199860
rect 148198 199832 148226 199940
rect 148290 199912 148318 200008
rect 148272 199860 148278 199912
rect 148330 199860 148336 199912
rect 148382 199832 148410 200076
rect 148658 200008 149330 200036
rect 148658 199912 148686 200008
rect 148548 199860 148554 199912
rect 148606 199860 148612 199912
rect 148640 199860 148646 199912
rect 148698 199860 148704 199912
rect 148916 199860 148922 199912
rect 148974 199860 148980 199912
rect 149100 199860 149106 199912
rect 149158 199860 149164 199912
rect 148198 199804 148410 199832
rect 148456 199792 148462 199844
rect 148514 199792 148520 199844
rect 148226 199696 148232 199708
rect 148106 199668 148232 199696
rect 148226 199656 148232 199668
rect 148284 199656 148290 199708
rect 147830 199600 147864 199640
rect 147858 199588 147864 199600
rect 147916 199588 147922 199640
rect 148134 199588 148140 199640
rect 148192 199628 148198 199640
rect 148474 199628 148502 199792
rect 148192 199600 148502 199628
rect 148192 199588 148198 199600
rect 148042 199520 148048 199572
rect 148100 199560 148106 199572
rect 148566 199560 148594 199860
rect 148934 199776 148962 199860
rect 148824 199724 148830 199776
rect 148882 199724 148888 199776
rect 148934 199736 148968 199776
rect 148962 199724 148968 199736
rect 149020 199724 149026 199776
rect 148842 199572 148870 199724
rect 148100 199532 148594 199560
rect 148100 199520 148106 199532
rect 148778 199520 148784 199572
rect 148836 199532 148870 199572
rect 148836 199520 148842 199532
rect 147858 199452 147864 199504
rect 147916 199492 147922 199504
rect 149118 199492 149146 199860
rect 147916 199464 149146 199492
rect 147916 199452 147922 199464
rect 148870 199316 148876 199368
rect 148928 199356 148934 199368
rect 149302 199356 149330 200008
rect 149376 199860 149382 199912
rect 149434 199900 149440 199912
rect 149434 199860 149468 199900
rect 149440 199776 149468 199860
rect 149422 199724 149428 199776
rect 149480 199724 149486 199776
rect 148928 199328 149330 199356
rect 148928 199316 148934 199328
rect 146628 199260 147628 199288
rect 149716 199288 149744 200416
rect 149836 199900 149842 199912
rect 149808 199860 149842 199900
rect 149894 199860 149900 199912
rect 150020 199860 150026 199912
rect 150078 199860 150084 199912
rect 150112 199860 150118 199912
rect 150170 199860 150176 199912
rect 150204 199860 150210 199912
rect 150262 199860 150268 199912
rect 150388 199860 150394 199912
rect 150446 199860 150452 199912
rect 150572 199860 150578 199912
rect 150630 199860 150636 199912
rect 149808 199504 149836 199860
rect 150038 199832 150066 199860
rect 149992 199804 150066 199832
rect 149992 199640 150020 199804
rect 150130 199776 150158 199860
rect 150066 199724 150072 199776
rect 150124 199736 150158 199776
rect 150124 199724 150130 199736
rect 150222 199708 150250 199860
rect 150406 199776 150434 199860
rect 150342 199724 150348 199776
rect 150400 199736 150434 199776
rect 150590 199776 150618 199860
rect 150774 199844 150802 200484
rect 151878 200348 153194 200376
rect 151004 200008 151630 200036
rect 150848 199860 150854 199912
rect 150906 199860 150912 199912
rect 150756 199792 150762 199844
rect 150814 199792 150820 199844
rect 150590 199736 150624 199776
rect 150400 199724 150406 199736
rect 150618 199724 150624 199736
rect 150676 199724 150682 199776
rect 150158 199656 150164 199708
rect 150216 199668 150250 199708
rect 150216 199656 150222 199668
rect 149974 199588 149980 199640
rect 150032 199588 150038 199640
rect 150250 199520 150256 199572
rect 150308 199560 150314 199572
rect 150710 199560 150716 199572
rect 150308 199532 150716 199560
rect 150308 199520 150314 199532
rect 150710 199520 150716 199532
rect 150768 199520 150774 199572
rect 149790 199452 149796 199504
rect 149848 199452 149854 199504
rect 150866 199356 150894 199860
rect 151004 199504 151032 200008
rect 151602 199968 151630 200008
rect 151602 199940 151722 199968
rect 151308 199900 151314 199912
rect 151280 199860 151314 199900
rect 151366 199860 151372 199912
rect 151400 199860 151406 199912
rect 151458 199860 151464 199912
rect 151584 199860 151590 199912
rect 151642 199860 151648 199912
rect 151124 199724 151130 199776
rect 151182 199724 151188 199776
rect 151142 199504 151170 199724
rect 151280 199696 151308 199860
rect 151418 199776 151446 199860
rect 151354 199724 151360 199776
rect 151412 199736 151446 199776
rect 151602 199764 151630 199860
rect 151694 199844 151722 199940
rect 151676 199792 151682 199844
rect 151734 199792 151740 199844
rect 151602 199736 151768 199764
rect 151412 199724 151418 199736
rect 151630 199696 151636 199708
rect 151280 199668 151636 199696
rect 151630 199656 151636 199668
rect 151688 199656 151694 199708
rect 151538 199520 151544 199572
rect 151596 199560 151602 199572
rect 151740 199560 151768 199736
rect 151596 199532 151768 199560
rect 151596 199520 151602 199532
rect 150986 199452 150992 199504
rect 151044 199452 151050 199504
rect 151142 199464 151176 199504
rect 151170 199452 151176 199464
rect 151228 199452 151234 199504
rect 151262 199452 151268 199504
rect 151320 199492 151326 199504
rect 151722 199492 151728 199504
rect 151320 199464 151728 199492
rect 151320 199452 151326 199464
rect 151722 199452 151728 199464
rect 151780 199452 151786 199504
rect 151630 199356 151636 199368
rect 150038 199328 150756 199356
rect 150866 199328 151636 199356
rect 150038 199288 150066 199328
rect 149716 199260 150066 199288
rect 146628 199248 146634 199260
rect 150250 199220 150256 199232
rect 145760 199192 150256 199220
rect 150250 199180 150256 199192
rect 150308 199180 150314 199232
rect 150434 199180 150440 199232
rect 150492 199220 150498 199232
rect 150728 199220 150756 199328
rect 151630 199316 151636 199328
rect 151688 199316 151694 199368
rect 150802 199248 150808 199300
rect 150860 199288 150866 199300
rect 151878 199288 151906 200348
rect 153166 200308 153194 200348
rect 159284 200308 159312 200552
rect 160066 200512 160094 200552
rect 161538 200512 161566 200688
rect 160066 200484 161106 200512
rect 161538 200484 161658 200512
rect 153166 200280 159312 200308
rect 150860 199260 151906 199288
rect 151970 200144 160922 200172
rect 150860 199248 150866 199260
rect 151970 199220 151998 200144
rect 152292 200008 154390 200036
rect 152292 199844 152320 200008
rect 153166 199940 153608 199968
rect 153166 199912 153194 199940
rect 152412 199860 152418 199912
rect 152470 199860 152476 199912
rect 153148 199860 153154 199912
rect 153206 199860 153212 199912
rect 153240 199860 153246 199912
rect 153298 199860 153304 199912
rect 152044 199792 152050 199844
rect 152102 199792 152108 199844
rect 152228 199792 152234 199844
rect 152286 199804 152320 199844
rect 152286 199792 152292 199804
rect 152062 199640 152090 199792
rect 152430 199696 152458 199860
rect 152596 199792 152602 199844
rect 152654 199792 152660 199844
rect 152780 199832 152786 199844
rect 152706 199804 152786 199832
rect 152384 199668 152458 199696
rect 152062 199600 152096 199640
rect 152090 199588 152096 199600
rect 152148 199588 152154 199640
rect 152384 199504 152412 199668
rect 152458 199588 152464 199640
rect 152516 199628 152522 199640
rect 152614 199628 152642 199792
rect 152516 199600 152642 199628
rect 152516 199588 152522 199600
rect 152366 199452 152372 199504
rect 152424 199452 152430 199504
rect 152706 199220 152734 199804
rect 152780 199792 152786 199804
rect 152838 199792 152844 199844
rect 152918 199696 152924 199708
rect 152844 199668 152924 199696
rect 152844 199640 152872 199668
rect 152918 199656 152924 199668
rect 152976 199656 152982 199708
rect 152826 199588 152832 199640
rect 152884 199588 152890 199640
rect 153258 199560 153286 199860
rect 153470 199560 153476 199572
rect 153258 199532 153476 199560
rect 153470 199520 153476 199532
rect 153528 199520 153534 199572
rect 153580 199492 153608 199940
rect 153212 199464 153608 199492
rect 153764 199940 154022 199968
rect 153764 199492 153792 199940
rect 153994 199912 154022 199940
rect 153884 199900 153890 199912
rect 153856 199860 153890 199900
rect 153942 199860 153948 199912
rect 153976 199860 153982 199912
rect 154034 199860 154040 199912
rect 154068 199860 154074 199912
rect 154126 199860 154132 199912
rect 154252 199860 154258 199912
rect 154310 199860 154316 199912
rect 153856 199696 153884 199860
rect 154086 199776 154114 199860
rect 154022 199724 154028 199776
rect 154080 199736 154114 199776
rect 154080 199724 154086 199736
rect 153856 199668 153976 199696
rect 153764 199464 153884 199492
rect 153212 199436 153240 199464
rect 153856 199436 153884 199464
rect 153194 199384 153200 199436
rect 153252 199384 153258 199436
rect 153378 199384 153384 199436
rect 153436 199424 153442 199436
rect 153746 199424 153752 199436
rect 153436 199396 153752 199424
rect 153436 199384 153442 199396
rect 153746 199384 153752 199396
rect 153804 199384 153810 199436
rect 153838 199384 153844 199436
rect 153896 199384 153902 199436
rect 150492 199180 150526 199220
rect 150728 199192 151998 199220
rect 152292 199192 152734 199220
rect 120258 199112 120264 199164
rect 120316 199152 120322 199164
rect 150498 199152 150526 199180
rect 151906 199152 151912 199164
rect 120316 199124 150434 199152
rect 150498 199124 151912 199152
rect 120316 199112 120322 199124
rect 125686 199044 125692 199096
rect 125744 199084 125750 199096
rect 135990 199084 135996 199096
rect 125744 199056 135996 199084
rect 125744 199044 125750 199056
rect 135990 199044 135996 199056
rect 136048 199044 136054 199096
rect 138934 199044 138940 199096
rect 138992 199084 138998 199096
rect 142982 199084 142988 199096
rect 138992 199056 142988 199084
rect 138992 199044 138998 199056
rect 142982 199044 142988 199056
rect 143040 199044 143046 199096
rect 145190 199044 145196 199096
rect 145248 199084 145254 199096
rect 150250 199084 150256 199096
rect 145248 199056 150256 199084
rect 145248 199044 145254 199056
rect 150250 199044 150256 199056
rect 150308 199044 150314 199096
rect 150406 199084 150434 199124
rect 151906 199112 151912 199124
rect 151964 199112 151970 199164
rect 152292 199084 152320 199192
rect 153102 199180 153108 199232
rect 153160 199220 153166 199232
rect 153948 199220 153976 199668
rect 154270 199640 154298 199860
rect 154206 199588 154212 199640
rect 154264 199600 154298 199640
rect 154362 199640 154390 200008
rect 158134 200008 160140 200036
rect 156294 199940 157656 199968
rect 156294 199912 156322 199940
rect 154436 199860 154442 199912
rect 154494 199860 154500 199912
rect 154620 199900 154626 199912
rect 154592 199860 154626 199900
rect 154678 199860 154684 199912
rect 154712 199860 154718 199912
rect 154770 199860 154776 199912
rect 154804 199860 154810 199912
rect 154862 199860 154868 199912
rect 154896 199860 154902 199912
rect 154954 199860 154960 199912
rect 154988 199860 154994 199912
rect 155046 199860 155052 199912
rect 155356 199860 155362 199912
rect 155414 199900 155420 199912
rect 155632 199900 155638 199912
rect 155414 199872 155540 199900
rect 155414 199860 155420 199872
rect 154454 199708 154482 199860
rect 154592 199708 154620 199860
rect 154730 199832 154758 199860
rect 154684 199804 154758 199832
rect 154684 199708 154712 199804
rect 154822 199764 154850 199860
rect 154776 199736 154850 199764
rect 154776 199708 154804 199736
rect 154914 199708 154942 199860
rect 154454 199668 154488 199708
rect 154482 199656 154488 199668
rect 154540 199656 154546 199708
rect 154574 199656 154580 199708
rect 154632 199656 154638 199708
rect 154666 199656 154672 199708
rect 154724 199656 154730 199708
rect 154758 199656 154764 199708
rect 154816 199656 154822 199708
rect 154850 199656 154856 199708
rect 154908 199668 154942 199708
rect 154908 199656 154914 199668
rect 154362 199600 154396 199640
rect 154264 199588 154270 199600
rect 154390 199588 154396 199600
rect 154448 199588 154454 199640
rect 155006 199560 155034 199860
rect 155512 199640 155540 199872
rect 155604 199860 155638 199900
rect 155690 199860 155696 199912
rect 155724 199860 155730 199912
rect 155782 199860 155788 199912
rect 156092 199860 156098 199912
rect 156150 199860 156156 199912
rect 156184 199860 156190 199912
rect 156242 199860 156248 199912
rect 156276 199860 156282 199912
rect 156334 199860 156340 199912
rect 156368 199860 156374 199912
rect 156426 199860 156432 199912
rect 156644 199900 156650 199912
rect 156524 199872 156650 199900
rect 155494 199588 155500 199640
rect 155552 199588 155558 199640
rect 155604 199628 155632 199860
rect 155742 199776 155770 199860
rect 155678 199724 155684 199776
rect 155736 199736 155770 199776
rect 155736 199724 155742 199736
rect 156110 199640 156138 199860
rect 156202 199708 156230 199860
rect 156386 199708 156414 199860
rect 156202 199668 156236 199708
rect 156230 199656 156236 199668
rect 156288 199656 156294 199708
rect 156322 199656 156328 199708
rect 156380 199668 156414 199708
rect 156380 199656 156386 199668
rect 156524 199640 156552 199872
rect 156644 199860 156650 199872
rect 156702 199860 156708 199912
rect 156736 199860 156742 199912
rect 156794 199860 156800 199912
rect 156828 199860 156834 199912
rect 156886 199860 156892 199912
rect 157104 199860 157110 199912
rect 157162 199900 157168 199912
rect 157162 199860 157196 199900
rect 157380 199860 157386 199912
rect 157438 199860 157444 199912
rect 156754 199832 156782 199860
rect 156616 199804 156782 199832
rect 155954 199628 155960 199640
rect 155604 199600 155960 199628
rect 155954 199588 155960 199600
rect 156012 199588 156018 199640
rect 156110 199600 156144 199640
rect 156138 199588 156144 199600
rect 156196 199588 156202 199640
rect 156506 199588 156512 199640
rect 156564 199588 156570 199640
rect 156616 199628 156644 199804
rect 156846 199776 156874 199860
rect 156920 199792 156926 199844
rect 156978 199792 156984 199844
rect 156782 199724 156788 199776
rect 156840 199736 156874 199776
rect 156840 199724 156846 199736
rect 156938 199640 156966 199792
rect 157058 199656 157064 199708
rect 157116 199696 157122 199708
rect 157168 199696 157196 199860
rect 157116 199668 157196 199696
rect 157116 199656 157122 199668
rect 157398 199640 157426 199860
rect 156690 199628 156696 199640
rect 156616 199600 156696 199628
rect 156690 199588 156696 199600
rect 156748 199588 156754 199640
rect 156938 199600 156972 199640
rect 156966 199588 156972 199600
rect 157024 199588 157030 199640
rect 157334 199588 157340 199640
rect 157392 199600 157426 199640
rect 157392 199588 157398 199600
rect 157628 199572 157656 199940
rect 158134 199912 158162 200008
rect 158272 199940 159542 199968
rect 157748 199860 157754 199912
rect 157806 199860 157812 199912
rect 157932 199900 157938 199912
rect 157904 199860 157938 199900
rect 157990 199860 157996 199912
rect 158024 199860 158030 199912
rect 158082 199860 158088 199912
rect 158116 199860 158122 199912
rect 158174 199860 158180 199912
rect 157766 199572 157794 199860
rect 157904 199572 157932 199860
rect 158042 199640 158070 199860
rect 158042 199600 158076 199640
rect 158070 199588 158076 199600
rect 158128 199588 158134 199640
rect 156874 199560 156880 199572
rect 155006 199532 156880 199560
rect 156874 199520 156880 199532
rect 156932 199520 156938 199572
rect 157610 199520 157616 199572
rect 157668 199520 157674 199572
rect 157702 199520 157708 199572
rect 157760 199532 157794 199572
rect 157760 199520 157766 199532
rect 157886 199520 157892 199572
rect 157944 199520 157950 199572
rect 155218 199452 155224 199504
rect 155276 199492 155282 199504
rect 158272 199492 158300 199940
rect 159514 199912 159542 199940
rect 158392 199900 158398 199912
rect 158364 199860 158398 199900
rect 158450 199860 158456 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158668 199860 158674 199912
rect 158726 199860 158732 199912
rect 159496 199860 159502 199912
rect 159554 199860 159560 199912
rect 159772 199860 159778 199912
rect 159830 199860 159836 199912
rect 159864 199860 159870 199912
rect 159922 199860 159928 199912
rect 158364 199708 158392 199860
rect 158502 199708 158530 199860
rect 158346 199656 158352 199708
rect 158404 199656 158410 199708
rect 158438 199656 158444 199708
rect 158496 199668 158530 199708
rect 158686 199696 158714 199860
rect 159790 199832 159818 199860
rect 158640 199668 158714 199696
rect 158962 199804 159818 199832
rect 158496 199656 158502 199668
rect 158640 199640 158668 199668
rect 158622 199588 158628 199640
rect 158680 199588 158686 199640
rect 158530 199520 158536 199572
rect 158588 199560 158594 199572
rect 158962 199560 158990 199804
rect 159882 199708 159910 199860
rect 159818 199656 159824 199708
rect 159876 199668 159910 199708
rect 159876 199656 159882 199668
rect 160112 199640 160140 200008
rect 160508 199900 160514 199912
rect 160204 199872 160514 199900
rect 160094 199588 160100 199640
rect 160152 199588 160158 199640
rect 158588 199532 158990 199560
rect 158588 199520 158594 199532
rect 158806 199492 158812 199504
rect 155276 199464 157288 199492
rect 158272 199464 158812 199492
rect 155276 199452 155282 199464
rect 156230 199384 156236 199436
rect 156288 199424 156294 199436
rect 157150 199424 157156 199436
rect 156288 199396 157156 199424
rect 156288 199384 156294 199396
rect 157150 199384 157156 199396
rect 157208 199384 157214 199436
rect 157260 199424 157288 199464
rect 158806 199452 158812 199464
rect 158864 199452 158870 199504
rect 160204 199492 160232 199872
rect 160508 199860 160514 199872
rect 160566 199860 160572 199912
rect 160692 199860 160698 199912
rect 160750 199860 160756 199912
rect 160784 199860 160790 199912
rect 160842 199860 160848 199912
rect 160324 199832 160330 199844
rect 160296 199792 160330 199832
rect 160382 199792 160388 199844
rect 160296 199708 160324 199792
rect 160416 199724 160422 199776
rect 160474 199724 160480 199776
rect 160710 199764 160738 199860
rect 160526 199736 160738 199764
rect 160278 199656 160284 199708
rect 160336 199656 160342 199708
rect 160434 199640 160462 199724
rect 160370 199588 160376 199640
rect 160428 199600 160462 199640
rect 160428 199588 160434 199600
rect 160526 199572 160554 199736
rect 160802 199696 160830 199860
rect 160462 199520 160468 199572
rect 160520 199532 160554 199572
rect 160756 199668 160830 199696
rect 160520 199520 160526 199532
rect 160066 199464 160232 199492
rect 160066 199424 160094 199464
rect 160554 199452 160560 199504
rect 160612 199492 160618 199504
rect 160756 199492 160784 199668
rect 160894 199640 160922 200144
rect 160968 199860 160974 199912
rect 161026 199860 161032 199912
rect 160830 199588 160836 199640
rect 160888 199600 160922 199640
rect 160888 199588 160894 199600
rect 160986 199572 161014 199860
rect 161078 199628 161106 200484
rect 161630 199912 161658 200484
rect 167334 200280 167776 200308
rect 163884 200008 164878 200036
rect 162780 199940 163314 199968
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161336 199860 161342 199912
rect 161394 199860 161400 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 161520 199860 161526 199912
rect 161578 199860 161584 199912
rect 161612 199860 161618 199912
rect 161670 199860 161676 199912
rect 161704 199860 161710 199912
rect 161762 199900 161768 199912
rect 161762 199860 161796 199900
rect 161888 199860 161894 199912
rect 161946 199860 161952 199912
rect 161980 199860 161986 199912
rect 162038 199860 162044 199912
rect 162072 199860 162078 199912
rect 162130 199860 162136 199912
rect 162256 199860 162262 199912
rect 162314 199900 162320 199912
rect 162314 199872 162716 199900
rect 162314 199860 162320 199872
rect 161170 199708 161198 199860
rect 161354 199776 161382 199860
rect 161290 199724 161296 199776
rect 161348 199736 161382 199776
rect 161348 199724 161354 199736
rect 161170 199668 161204 199708
rect 161198 199656 161204 199668
rect 161256 199656 161262 199708
rect 161446 199640 161474 199860
rect 161538 199776 161566 199860
rect 161630 199832 161658 199860
rect 161630 199804 161704 199832
rect 161538 199736 161572 199776
rect 161566 199724 161572 199736
rect 161624 199724 161630 199776
rect 161078 199600 161152 199628
rect 160986 199532 161020 199572
rect 161014 199520 161020 199532
rect 161072 199520 161078 199572
rect 161124 199492 161152 199600
rect 161382 199588 161388 199640
rect 161440 199600 161474 199640
rect 161440 199588 161446 199600
rect 160612 199464 160784 199492
rect 160986 199464 161152 199492
rect 160612 199452 160618 199464
rect 157260 199396 160094 199424
rect 160738 199384 160744 199436
rect 160796 199424 160802 199436
rect 160986 199424 161014 199464
rect 160796 199396 161014 199424
rect 160796 199384 160802 199396
rect 154942 199316 154948 199368
rect 155000 199356 155006 199368
rect 157334 199356 157340 199368
rect 155000 199328 157340 199356
rect 155000 199316 155006 199328
rect 157334 199316 157340 199328
rect 157392 199316 157398 199368
rect 161676 199356 161704 199804
rect 161768 199640 161796 199860
rect 161750 199588 161756 199640
rect 161808 199588 161814 199640
rect 161906 199560 161934 199860
rect 161998 199640 162026 199860
rect 162090 199696 162118 199860
rect 162090 199668 162440 199696
rect 161998 199600 162032 199640
rect 162026 199588 162032 199600
rect 162084 199588 162090 199640
rect 162412 199628 162440 199668
rect 162412 199600 162624 199628
rect 162486 199560 162492 199572
rect 161906 199532 162492 199560
rect 162486 199520 162492 199532
rect 162544 199520 162550 199572
rect 161934 199452 161940 199504
rect 161992 199492 161998 199504
rect 162596 199492 162624 199600
rect 161992 199464 162624 199492
rect 161992 199452 161998 199464
rect 162210 199384 162216 199436
rect 162268 199424 162274 199436
rect 162688 199424 162716 199872
rect 162780 199640 162808 199940
rect 163286 199912 163314 199940
rect 162900 199860 162906 199912
rect 162958 199860 162964 199912
rect 163084 199900 163090 199912
rect 163056 199860 163090 199900
rect 163142 199860 163148 199912
rect 163176 199860 163182 199912
rect 163234 199860 163240 199912
rect 163268 199860 163274 199912
rect 163326 199860 163332 199912
rect 163728 199860 163734 199912
rect 163786 199860 163792 199912
rect 162762 199588 162768 199640
rect 162820 199588 162826 199640
rect 162918 199492 162946 199860
rect 163056 199640 163084 199860
rect 163194 199832 163222 199860
rect 163148 199804 163222 199832
rect 163038 199588 163044 199640
rect 163096 199588 163102 199640
rect 163148 199560 163176 199804
rect 163746 199628 163774 199860
rect 163332 199600 163774 199628
rect 163222 199560 163228 199572
rect 163148 199532 163228 199560
rect 163222 199520 163228 199532
rect 163280 199520 163286 199572
rect 163038 199492 163044 199504
rect 162918 199464 163044 199492
rect 163038 199452 163044 199464
rect 163096 199452 163102 199504
rect 163332 199492 163360 199600
rect 163774 199492 163780 199504
rect 163332 199464 163780 199492
rect 163774 199452 163780 199464
rect 163832 199452 163838 199504
rect 162268 199396 162716 199424
rect 163884 199424 163912 200008
rect 164390 199940 164694 199968
rect 164188 199860 164194 199912
rect 164246 199860 164252 199912
rect 164096 199792 164102 199844
rect 164154 199792 164160 199844
rect 164114 199764 164142 199792
rect 164068 199736 164142 199764
rect 164068 199708 164096 199736
rect 164206 199708 164234 199860
rect 164050 199656 164056 199708
rect 164108 199656 164114 199708
rect 164142 199656 164148 199708
rect 164200 199668 164234 199708
rect 164200 199656 164206 199668
rect 163958 199452 163964 199504
rect 164016 199492 164022 199504
rect 164234 199492 164240 199504
rect 164016 199464 164240 199492
rect 164016 199452 164022 199464
rect 164234 199452 164240 199464
rect 164292 199452 164298 199504
rect 164390 199492 164418 199940
rect 164666 199912 164694 199940
rect 164850 199912 164878 200008
rect 165264 200008 166074 200036
rect 164464 199860 164470 199912
rect 164522 199860 164528 199912
rect 164648 199860 164654 199912
rect 164706 199860 164712 199912
rect 164740 199860 164746 199912
rect 164798 199860 164804 199912
rect 164832 199860 164838 199912
rect 164890 199860 164896 199912
rect 164924 199860 164930 199912
rect 164982 199860 164988 199912
rect 165108 199860 165114 199912
rect 165166 199860 165172 199912
rect 164482 199560 164510 199860
rect 164758 199696 164786 199860
rect 164942 199708 164970 199860
rect 164758 199668 164832 199696
rect 164694 199560 164700 199572
rect 164482 199532 164700 199560
rect 164694 199520 164700 199532
rect 164752 199520 164758 199572
rect 164510 199492 164516 199504
rect 164390 199464 164516 199492
rect 164510 199452 164516 199464
rect 164568 199452 164574 199504
rect 164602 199452 164608 199504
rect 164660 199492 164666 199504
rect 164804 199492 164832 199668
rect 164878 199656 164884 199708
rect 164936 199668 164970 199708
rect 164936 199656 164942 199668
rect 165126 199640 165154 199860
rect 165062 199588 165068 199640
rect 165120 199600 165154 199640
rect 165120 199588 165126 199600
rect 164660 199464 164832 199492
rect 164660 199452 164666 199464
rect 164878 199452 164884 199504
rect 164936 199492 164942 199504
rect 165264 199492 165292 200008
rect 165844 199860 165850 199912
rect 165902 199860 165908 199912
rect 165936 199860 165942 199912
rect 165994 199900 166000 199912
rect 166046 199900 166074 200008
rect 166414 199940 166718 199968
rect 165994 199872 166074 199900
rect 165994 199860 166000 199872
rect 166120 199860 166126 199912
rect 166178 199860 166184 199912
rect 165862 199696 165890 199860
rect 166138 199832 166166 199860
rect 166092 199804 166166 199832
rect 166092 199776 166120 199804
rect 166304 199792 166310 199844
rect 166362 199792 166368 199844
rect 166074 199724 166080 199776
rect 166132 199724 166138 199776
rect 166322 199708 166350 199792
rect 165982 199696 165988 199708
rect 165862 199668 165988 199696
rect 165982 199656 165988 199668
rect 166040 199656 166046 199708
rect 166258 199656 166264 199708
rect 166316 199668 166350 199708
rect 166316 199656 166322 199668
rect 166414 199560 166442 199940
rect 166690 199912 166718 199940
rect 166672 199860 166678 199912
rect 166730 199860 166736 199912
rect 166764 199860 166770 199912
rect 166822 199860 166828 199912
rect 167132 199860 167138 199912
rect 167190 199860 167196 199912
rect 167224 199860 167230 199912
rect 167282 199860 167288 199912
rect 166782 199776 166810 199860
rect 167040 199832 167046 199844
rect 166718 199724 166724 199776
rect 166776 199736 166810 199776
rect 166874 199804 167046 199832
rect 166776 199724 166782 199736
rect 166874 199696 166902 199804
rect 167040 199792 167046 199804
rect 167098 199792 167104 199844
rect 167150 199708 167178 199860
rect 164936 199464 165292 199492
rect 165816 199532 166442 199560
rect 166690 199668 166902 199696
rect 164936 199452 164942 199464
rect 165246 199424 165252 199436
rect 163884 199396 165252 199424
rect 162268 199384 162274 199396
rect 165246 199384 165252 199396
rect 165304 199384 165310 199436
rect 165430 199356 165436 199368
rect 161676 199328 165436 199356
rect 165430 199316 165436 199328
rect 165488 199316 165494 199368
rect 165816 199356 165844 199532
rect 165890 199384 165896 199436
rect 165948 199424 165954 199436
rect 166690 199424 166718 199668
rect 167086 199656 167092 199708
rect 167144 199668 167178 199708
rect 167144 199656 167150 199668
rect 167242 199628 167270 199860
rect 165948 199396 166718 199424
rect 166920 199600 167270 199628
rect 165948 199384 165954 199396
rect 166626 199356 166632 199368
rect 165816 199328 166632 199356
rect 166626 199316 166632 199328
rect 166684 199316 166690 199368
rect 166920 199356 166948 199600
rect 167334 199572 167362 200280
rect 167748 199912 167776 200280
rect 167840 199968 167868 200756
rect 169358 200756 580724 200784
rect 169358 199968 169386 200756
rect 580718 200744 580724 200756
rect 580776 200744 580782 200796
rect 562318 200716 562324 200728
rect 171106 200688 562324 200716
rect 171106 200580 171134 200688
rect 562318 200676 562324 200688
rect 562376 200676 562382 200728
rect 177942 200608 177948 200660
rect 178000 200648 178006 200660
rect 191742 200648 191748 200660
rect 178000 200620 191748 200648
rect 178000 200608 178006 200620
rect 191742 200608 191748 200620
rect 191800 200608 191806 200660
rect 169726 200552 171134 200580
rect 179386 200552 182174 200580
rect 167840 199940 169110 199968
rect 169358 199940 169478 199968
rect 167408 199860 167414 199912
rect 167466 199860 167472 199912
rect 167748 199872 167782 199912
rect 167776 199860 167782 199872
rect 167834 199860 167840 199912
rect 167868 199860 167874 199912
rect 167926 199860 167932 199912
rect 167960 199860 167966 199912
rect 168018 199860 168024 199912
rect 168052 199860 168058 199912
rect 168110 199860 168116 199912
rect 168144 199860 168150 199912
rect 168202 199900 168208 199912
rect 168202 199860 168236 199900
rect 168328 199860 168334 199912
rect 168386 199860 168392 199912
rect 168420 199860 168426 199912
rect 168478 199860 168484 199912
rect 167270 199520 167276 199572
rect 167328 199532 167362 199572
rect 167328 199520 167334 199532
rect 167426 199492 167454 199860
rect 167638 199520 167644 199572
rect 167696 199560 167702 199572
rect 167886 199560 167914 199860
rect 167696 199532 167914 199560
rect 167978 199572 168006 199860
rect 168070 199628 168098 199860
rect 168070 199600 168144 199628
rect 168116 199572 168144 199600
rect 167978 199532 168012 199572
rect 167696 199520 167702 199532
rect 168006 199520 168012 199532
rect 168064 199520 168070 199572
rect 168098 199520 168104 199572
rect 168156 199520 168162 199572
rect 167914 199492 167920 199504
rect 167426 199464 167920 199492
rect 167914 199452 167920 199464
rect 167972 199452 167978 199504
rect 167178 199384 167184 199436
rect 167236 199424 167242 199436
rect 168208 199424 168236 199860
rect 168346 199832 168374 199860
rect 167236 199396 168236 199424
rect 168300 199804 168374 199832
rect 168300 199424 168328 199804
rect 168438 199708 168466 199860
rect 168374 199656 168380 199708
rect 168432 199668 168466 199708
rect 168432 199656 168438 199668
rect 168576 199640 168604 199940
rect 169082 199912 169110 199940
rect 169064 199860 169070 199912
rect 169122 199860 169128 199912
rect 169340 199860 169346 199912
rect 169398 199860 169404 199912
rect 169358 199776 169386 199860
rect 169294 199724 169300 199776
rect 169352 199736 169386 199776
rect 169352 199724 169358 199736
rect 168558 199588 168564 199640
rect 168616 199588 168622 199640
rect 169110 199588 169116 199640
rect 169168 199628 169174 199640
rect 169450 199628 169478 199940
rect 169616 199860 169622 199912
rect 169674 199860 169680 199912
rect 169634 199708 169662 199860
rect 169616 199656 169622 199708
rect 169674 199656 169680 199708
rect 169168 199600 169478 199628
rect 169168 199588 169174 199600
rect 169386 199520 169392 199572
rect 169444 199560 169450 199572
rect 169726 199560 169754 200552
rect 179386 200512 179414 200552
rect 169818 200484 179414 200512
rect 169818 199912 169846 200484
rect 178678 200444 178684 200456
rect 173866 200416 178684 200444
rect 171382 199940 172100 199968
rect 171382 199912 171410 199940
rect 169800 199860 169806 199912
rect 169858 199860 169864 199912
rect 169984 199900 169990 199912
rect 169956 199860 169990 199900
rect 170042 199860 170048 199912
rect 170076 199860 170082 199912
rect 170134 199860 170140 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 170444 199860 170450 199912
rect 170502 199860 170508 199912
rect 170536 199860 170542 199912
rect 170594 199860 170600 199912
rect 170996 199860 171002 199912
rect 171054 199860 171060 199912
rect 171272 199860 171278 199912
rect 171330 199860 171336 199912
rect 171364 199860 171370 199912
rect 171422 199860 171428 199912
rect 171456 199860 171462 199912
rect 171514 199860 171520 199912
rect 171824 199860 171830 199912
rect 171882 199860 171888 199912
rect 171916 199860 171922 199912
rect 171974 199900 171980 199912
rect 171974 199860 172008 199900
rect 169956 199776 169984 199860
rect 170094 199832 170122 199860
rect 170048 199804 170122 199832
rect 169938 199724 169944 199776
rect 169996 199724 170002 199776
rect 170048 199708 170076 199804
rect 170186 199776 170214 199860
rect 170122 199724 170128 199776
rect 170180 199736 170214 199776
rect 170462 199776 170490 199860
rect 170554 199832 170582 199860
rect 170554 199804 170628 199832
rect 170600 199776 170628 199804
rect 171014 199776 171042 199860
rect 170462 199736 170496 199776
rect 170180 199724 170186 199736
rect 170490 199724 170496 199736
rect 170548 199724 170554 199776
rect 170582 199724 170588 199776
rect 170640 199724 170646 199776
rect 170950 199724 170956 199776
rect 171008 199736 171042 199776
rect 171008 199724 171014 199736
rect 170030 199656 170036 199708
rect 170088 199656 170094 199708
rect 171290 199696 171318 199860
rect 171474 199776 171502 199860
rect 171410 199724 171416 199776
rect 171468 199736 171502 199776
rect 171468 199724 171474 199736
rect 171152 199668 171318 199696
rect 169444 199532 169754 199560
rect 171152 199560 171180 199668
rect 171594 199560 171600 199572
rect 171152 199532 171600 199560
rect 169444 199520 169450 199532
rect 171594 199520 171600 199532
rect 171652 199520 171658 199572
rect 171842 199560 171870 199860
rect 171980 199776 172008 199860
rect 171962 199724 171968 199776
rect 172020 199724 172026 199776
rect 171704 199532 171870 199560
rect 172072 199560 172100 199940
rect 172376 199860 172382 199912
rect 172434 199860 172440 199912
rect 172560 199860 172566 199912
rect 172618 199900 172624 199912
rect 172618 199860 172652 199900
rect 172836 199860 172842 199912
rect 172894 199860 172900 199912
rect 172928 199860 172934 199912
rect 172986 199860 172992 199912
rect 173020 199860 173026 199912
rect 173078 199860 173084 199912
rect 173204 199860 173210 199912
rect 173262 199860 173268 199912
rect 173480 199860 173486 199912
rect 173538 199860 173544 199912
rect 173664 199860 173670 199912
rect 173722 199900 173728 199912
rect 173866 199900 173894 200416
rect 178678 200404 178684 200416
rect 178736 200404 178742 200456
rect 182146 200308 182174 200552
rect 182146 200280 183554 200308
rect 178770 200240 178776 200252
rect 173958 200212 178776 200240
rect 173958 199912 173986 200212
rect 178770 200200 178776 200212
rect 178828 200200 178834 200252
rect 183526 200172 183554 200280
rect 194502 200268 194508 200320
rect 194560 200308 194566 200320
rect 211430 200308 211436 200320
rect 194560 200280 211436 200308
rect 194560 200268 194566 200280
rect 211430 200268 211436 200280
rect 211488 200268 211494 200320
rect 190546 200200 190552 200252
rect 190604 200240 190610 200252
rect 191650 200240 191656 200252
rect 190604 200212 191656 200240
rect 190604 200200 190610 200212
rect 191650 200200 191656 200212
rect 191708 200240 191714 200252
rect 215386 200240 215392 200252
rect 191708 200212 215392 200240
rect 191708 200200 191714 200212
rect 215386 200200 215392 200212
rect 215444 200200 215450 200252
rect 204346 200172 204352 200184
rect 183526 200144 204352 200172
rect 204346 200132 204352 200144
rect 204404 200132 204410 200184
rect 178402 200104 178408 200116
rect 174602 200076 178408 200104
rect 174602 199912 174630 200076
rect 178402 200064 178408 200076
rect 178460 200064 178466 200116
rect 180518 200036 180524 200048
rect 175384 200008 180524 200036
rect 174878 199940 175090 199968
rect 173722 199872 173894 199900
rect 173722 199860 173728 199872
rect 173940 199860 173946 199912
rect 173998 199860 174004 199912
rect 174032 199860 174038 199912
rect 174090 199860 174096 199912
rect 174124 199860 174130 199912
rect 174182 199860 174188 199912
rect 174400 199860 174406 199912
rect 174458 199860 174464 199912
rect 174584 199860 174590 199912
rect 174642 199860 174648 199912
rect 174768 199860 174774 199912
rect 174826 199860 174832 199912
rect 172192 199724 172198 199776
rect 172250 199724 172256 199776
rect 172210 199640 172238 199724
rect 172394 199708 172422 199860
rect 172394 199668 172428 199708
rect 172422 199656 172428 199668
rect 172480 199656 172486 199708
rect 172624 199640 172652 199860
rect 172854 199776 172882 199860
rect 172790 199724 172796 199776
rect 172848 199736 172882 199776
rect 172848 199724 172854 199736
rect 172946 199708 172974 199860
rect 172882 199656 172888 199708
rect 172940 199668 172974 199708
rect 172940 199656 172946 199668
rect 173038 199640 173066 199860
rect 173222 199776 173250 199860
rect 173158 199724 173164 199776
rect 173216 199736 173250 199776
rect 173216 199724 173222 199736
rect 172146 199588 172152 199640
rect 172204 199600 172238 199640
rect 172204 199588 172210 199600
rect 172606 199588 172612 199640
rect 172664 199588 172670 199640
rect 172974 199588 172980 199640
rect 173032 199600 173066 199640
rect 173498 199640 173526 199860
rect 174050 199776 174078 199860
rect 173986 199724 173992 199776
rect 174044 199736 174078 199776
rect 174044 199724 174050 199736
rect 173848 199656 173854 199708
rect 173906 199656 173912 199708
rect 174142 199696 174170 199860
rect 174418 199832 174446 199860
rect 174418 199804 174492 199832
rect 174464 199776 174492 199804
rect 174786 199776 174814 199860
rect 174446 199724 174452 199776
rect 174504 199724 174510 199776
rect 174722 199724 174728 199776
rect 174780 199736 174814 199776
rect 174780 199724 174786 199736
rect 174630 199696 174636 199708
rect 174142 199668 174636 199696
rect 174630 199656 174636 199668
rect 174688 199656 174694 199708
rect 173498 199600 173532 199640
rect 173032 199588 173038 199600
rect 173526 199588 173532 199600
rect 173584 199588 173590 199640
rect 173866 199628 173894 199656
rect 173866 199600 174308 199628
rect 174280 199572 174308 199600
rect 174878 199572 174906 199940
rect 175062 199912 175090 199940
rect 175384 199912 175412 200008
rect 180518 199996 180524 200008
rect 180576 199996 180582 200048
rect 181806 199968 181812 199980
rect 176350 199940 176654 199968
rect 174952 199860 174958 199912
rect 175010 199860 175016 199912
rect 175044 199860 175050 199912
rect 175102 199860 175108 199912
rect 175136 199860 175142 199912
rect 175194 199860 175200 199912
rect 175228 199860 175234 199912
rect 175286 199860 175292 199912
rect 175384 199872 175418 199912
rect 175412 199860 175418 199872
rect 175470 199860 175476 199912
rect 175688 199900 175694 199912
rect 175660 199860 175694 199900
rect 175746 199860 175752 199912
rect 176148 199860 176154 199912
rect 176206 199860 176212 199912
rect 174970 199628 174998 199860
rect 175154 199776 175182 199860
rect 175090 199724 175096 199776
rect 175148 199736 175182 199776
rect 175148 199724 175154 199736
rect 175090 199628 175096 199640
rect 174970 199600 175096 199628
rect 175090 199588 175096 199600
rect 175148 199588 175154 199640
rect 172238 199560 172244 199572
rect 172072 199532 172244 199560
rect 168466 199452 168472 199504
rect 168524 199492 168530 199504
rect 169662 199492 169668 199504
rect 168524 199464 169668 199492
rect 168524 199452 168530 199464
rect 169662 199452 169668 199464
rect 169720 199452 169726 199504
rect 171226 199452 171232 199504
rect 171284 199492 171290 199504
rect 171704 199492 171732 199532
rect 172238 199520 172244 199532
rect 172296 199520 172302 199572
rect 174262 199520 174268 199572
rect 174320 199520 174326 199572
rect 174878 199532 174912 199572
rect 174906 199520 174912 199532
rect 174964 199520 174970 199572
rect 174998 199520 175004 199572
rect 175056 199560 175062 199572
rect 175246 199560 175274 199860
rect 175320 199724 175326 199776
rect 175378 199764 175384 199776
rect 175378 199724 175412 199764
rect 175384 199640 175412 199724
rect 175366 199588 175372 199640
rect 175424 199588 175430 199640
rect 175660 199628 175688 199860
rect 175872 199832 175878 199844
rect 175752 199804 175878 199832
rect 175752 199708 175780 199804
rect 175872 199792 175878 199804
rect 175930 199792 175936 199844
rect 175734 199656 175740 199708
rect 175792 199656 175798 199708
rect 175826 199656 175832 199708
rect 175884 199696 175890 199708
rect 176166 199696 176194 199860
rect 176350 199844 176378 199940
rect 176516 199860 176522 199912
rect 176574 199860 176580 199912
rect 176332 199792 176338 199844
rect 176390 199792 176396 199844
rect 175884 199668 176194 199696
rect 175884 199656 175890 199668
rect 176286 199628 176292 199640
rect 175660 199600 176292 199628
rect 176286 199588 176292 199600
rect 176344 199588 176350 199640
rect 176378 199588 176384 199640
rect 176436 199628 176442 199640
rect 176534 199628 176562 199860
rect 176626 199696 176654 199940
rect 177178 199940 181812 199968
rect 177178 199912 177206 199940
rect 181806 199928 181812 199940
rect 181864 199928 181870 199980
rect 176700 199860 176706 199912
rect 176758 199900 176764 199912
rect 176758 199872 177114 199900
rect 176758 199860 176764 199872
rect 177086 199832 177114 199872
rect 177160 199860 177166 199912
rect 177218 199860 177224 199912
rect 177344 199860 177350 199912
rect 177402 199900 177408 199912
rect 180426 199900 180432 199912
rect 177402 199872 180432 199900
rect 177402 199860 177408 199872
rect 180426 199860 180432 199872
rect 180484 199860 180490 199912
rect 178034 199832 178040 199844
rect 177086 199804 178040 199832
rect 178034 199792 178040 199804
rect 178092 199792 178098 199844
rect 177666 199724 177672 199776
rect 177724 199764 177730 199776
rect 188982 199764 188988 199776
rect 177724 199736 188988 199764
rect 177724 199724 177730 199736
rect 188982 199724 188988 199736
rect 189040 199764 189046 199776
rect 192478 199764 192484 199776
rect 189040 199736 192484 199764
rect 189040 199724 189046 199736
rect 192478 199724 192484 199736
rect 192536 199724 192542 199776
rect 182266 199696 182272 199708
rect 176626 199668 182272 199696
rect 182266 199656 182272 199668
rect 182324 199656 182330 199708
rect 176436 199600 176562 199628
rect 176436 199588 176442 199600
rect 178954 199588 178960 199640
rect 179012 199628 179018 199640
rect 302234 199628 302240 199640
rect 179012 199600 302240 199628
rect 179012 199588 179018 199600
rect 302234 199588 302240 199600
rect 302292 199588 302298 199640
rect 184750 199560 184756 199572
rect 175056 199532 175274 199560
rect 176120 199532 184756 199560
rect 175056 199520 175062 199532
rect 171284 199464 171732 199492
rect 171284 199452 171290 199464
rect 171778 199452 171784 199504
rect 171836 199492 171842 199504
rect 176120 199492 176148 199532
rect 184750 199520 184756 199532
rect 184808 199560 184814 199572
rect 189810 199560 189816 199572
rect 184808 199532 189816 199560
rect 184808 199520 184814 199532
rect 189810 199520 189816 199532
rect 189868 199520 189874 199572
rect 199378 199560 199384 199572
rect 190426 199532 199384 199560
rect 171836 199464 176148 199492
rect 171836 199452 171842 199464
rect 176654 199452 176660 199504
rect 176712 199492 176718 199504
rect 176930 199492 176936 199504
rect 176712 199464 176936 199492
rect 176712 199452 176718 199464
rect 176930 199452 176936 199464
rect 176988 199452 176994 199504
rect 184934 199452 184940 199504
rect 184992 199492 184998 199504
rect 186222 199492 186228 199504
rect 184992 199464 186228 199492
rect 184992 199452 184998 199464
rect 186222 199452 186228 199464
rect 186280 199492 186286 199504
rect 190426 199492 190454 199532
rect 199378 199520 199384 199532
rect 199436 199520 199442 199572
rect 216674 199520 216680 199572
rect 216732 199560 216738 199572
rect 427814 199560 427820 199572
rect 216732 199532 427820 199560
rect 216732 199520 216738 199532
rect 427814 199520 427820 199532
rect 427872 199520 427878 199572
rect 186280 199464 190454 199492
rect 186280 199452 186286 199464
rect 201402 199452 201408 199504
rect 201460 199492 201466 199504
rect 412634 199492 412640 199504
rect 201460 199464 412640 199492
rect 201460 199452 201466 199464
rect 412634 199452 412640 199464
rect 412692 199452 412698 199504
rect 168650 199424 168656 199436
rect 168300 199396 168656 199424
rect 167236 199384 167242 199396
rect 168650 199384 168656 199396
rect 168708 199384 168714 199436
rect 170766 199384 170772 199436
rect 170824 199424 170830 199436
rect 431954 199424 431960 199436
rect 170824 199396 431960 199424
rect 170824 199384 170830 199396
rect 431954 199384 431960 199396
rect 432012 199384 432018 199436
rect 167362 199356 167368 199368
rect 166920 199328 167368 199356
rect 167362 199316 167368 199328
rect 167420 199316 167426 199368
rect 170306 199316 170312 199368
rect 170364 199356 170370 199368
rect 182174 199356 182180 199368
rect 170364 199328 182180 199356
rect 170364 199316 170370 199328
rect 182174 199316 182180 199328
rect 182232 199316 182238 199368
rect 156230 199248 156236 199300
rect 156288 199288 156294 199300
rect 156966 199288 156972 199300
rect 156288 199260 156972 199288
rect 156288 199248 156294 199260
rect 156966 199248 156972 199260
rect 157024 199248 157030 199300
rect 157242 199248 157248 199300
rect 157300 199288 157306 199300
rect 291194 199288 291200 199300
rect 157300 199260 291200 199288
rect 157300 199248 157306 199260
rect 291194 199248 291200 199260
rect 291252 199248 291258 199300
rect 153160 199192 153976 199220
rect 153160 199180 153166 199192
rect 159634 199180 159640 199232
rect 159692 199220 159698 199232
rect 216674 199220 216680 199232
rect 159692 199192 216680 199220
rect 159692 199180 159698 199192
rect 216674 199180 216680 199192
rect 216732 199180 216738 199232
rect 152734 199112 152740 199164
rect 152792 199152 152798 199164
rect 154022 199152 154028 199164
rect 152792 199124 154028 199152
rect 152792 199112 152798 199124
rect 154022 199112 154028 199124
rect 154080 199112 154086 199164
rect 155494 199112 155500 199164
rect 155552 199152 155558 199164
rect 190546 199152 190552 199164
rect 155552 199124 190552 199152
rect 155552 199112 155558 199124
rect 190546 199112 190552 199124
rect 190604 199112 190610 199164
rect 150406 199056 152320 199084
rect 152642 199044 152648 199096
rect 152700 199084 152706 199096
rect 154942 199084 154948 199096
rect 152700 199056 154948 199084
rect 152700 199044 152706 199056
rect 154942 199044 154948 199056
rect 155000 199044 155006 199096
rect 160094 199044 160100 199096
rect 160152 199084 160158 199096
rect 184934 199084 184940 199096
rect 160152 199056 184940 199084
rect 160152 199044 160158 199056
rect 184934 199044 184940 199056
rect 184992 199044 184998 199096
rect 130378 198976 130384 199028
rect 130436 199016 130442 199028
rect 147950 199016 147956 199028
rect 130436 198988 147956 199016
rect 130436 198976 130442 198988
rect 147950 198976 147956 198988
rect 148008 199016 148014 199028
rect 190086 199016 190092 199028
rect 148008 198988 190092 199016
rect 148008 198976 148014 198988
rect 190086 198976 190092 198988
rect 190144 198976 190150 199028
rect 117958 198908 117964 198960
rect 118016 198948 118022 198960
rect 164050 198948 164056 198960
rect 118016 198920 164056 198948
rect 118016 198908 118022 198920
rect 164050 198908 164056 198920
rect 164108 198908 164114 198960
rect 164234 198908 164240 198960
rect 164292 198948 164298 198960
rect 164786 198948 164792 198960
rect 164292 198920 164792 198948
rect 164292 198908 164298 198920
rect 164786 198908 164792 198920
rect 164844 198908 164850 198960
rect 175550 198948 175556 198960
rect 164896 198920 175556 198948
rect 120718 198840 120724 198892
rect 120776 198880 120782 198892
rect 124306 198880 124312 198892
rect 120776 198852 124312 198880
rect 120776 198840 120782 198852
rect 124306 198840 124312 198852
rect 124364 198880 124370 198892
rect 125502 198880 125508 198892
rect 124364 198852 125508 198880
rect 124364 198840 124370 198852
rect 125502 198840 125508 198852
rect 125560 198840 125566 198892
rect 128906 198840 128912 198892
rect 128964 198880 128970 198892
rect 133138 198880 133144 198892
rect 128964 198852 133144 198880
rect 128964 198840 128970 198852
rect 133138 198840 133144 198852
rect 133196 198840 133202 198892
rect 135898 198840 135904 198892
rect 135956 198880 135962 198892
rect 140958 198880 140964 198892
rect 135956 198852 140964 198880
rect 135956 198840 135962 198852
rect 140958 198840 140964 198852
rect 141016 198840 141022 198892
rect 142706 198840 142712 198892
rect 142764 198880 142770 198892
rect 145190 198880 145196 198892
rect 142764 198852 145196 198880
rect 142764 198840 142770 198852
rect 145190 198840 145196 198852
rect 145248 198840 145254 198892
rect 145650 198840 145656 198892
rect 145708 198880 145714 198892
rect 157242 198880 157248 198892
rect 145708 198852 157248 198880
rect 145708 198840 145714 198852
rect 157242 198840 157248 198852
rect 157300 198840 157306 198892
rect 160830 198840 160836 198892
rect 160888 198880 160894 198892
rect 163590 198880 163596 198892
rect 160888 198852 163596 198880
rect 160888 198840 160894 198852
rect 163590 198840 163596 198852
rect 163648 198840 163654 198892
rect 120902 198772 120908 198824
rect 120960 198812 120966 198824
rect 164896 198812 164924 198920
rect 175550 198908 175556 198920
rect 175608 198948 175614 198960
rect 175826 198948 175832 198960
rect 175608 198920 175832 198948
rect 175608 198908 175614 198920
rect 175826 198908 175832 198920
rect 175884 198908 175890 198960
rect 176194 198908 176200 198960
rect 176252 198948 176258 198960
rect 176562 198948 176568 198960
rect 176252 198920 176568 198948
rect 176252 198908 176258 198920
rect 176562 198908 176568 198920
rect 176620 198908 176626 198960
rect 178034 198908 178040 198960
rect 178092 198948 178098 198960
rect 178092 198920 182174 198948
rect 178092 198908 178098 198920
rect 165430 198840 165436 198892
rect 165488 198880 165494 198892
rect 166166 198880 166172 198892
rect 165488 198852 166172 198880
rect 165488 198840 165494 198852
rect 166166 198840 166172 198852
rect 166224 198840 166230 198892
rect 169202 198840 169208 198892
rect 169260 198880 169266 198892
rect 169260 198852 173894 198880
rect 169260 198840 169266 198852
rect 120960 198784 146616 198812
rect 120960 198772 120966 198784
rect 120810 198704 120816 198756
rect 120868 198744 120874 198756
rect 124766 198744 124772 198756
rect 120868 198716 124772 198744
rect 120868 198704 120874 198716
rect 124766 198704 124772 198716
rect 124824 198704 124830 198756
rect 125502 198704 125508 198756
rect 125560 198744 125566 198756
rect 144546 198744 144552 198756
rect 125560 198716 144552 198744
rect 125560 198704 125566 198716
rect 144546 198704 144552 198716
rect 144604 198704 144610 198756
rect 120718 198636 120724 198688
rect 120776 198676 120782 198688
rect 120776 198648 122834 198676
rect 120776 198636 120782 198648
rect 121178 198568 121184 198620
rect 121236 198608 121242 198620
rect 122806 198608 122834 198648
rect 126514 198636 126520 198688
rect 126572 198676 126578 198688
rect 134518 198676 134524 198688
rect 126572 198648 134524 198676
rect 126572 198636 126578 198648
rect 134518 198636 134524 198648
rect 134576 198636 134582 198688
rect 136266 198636 136272 198688
rect 136324 198676 136330 198688
rect 143994 198676 144000 198688
rect 136324 198648 144000 198676
rect 136324 198636 136330 198648
rect 143994 198636 144000 198648
rect 144052 198636 144058 198688
rect 138382 198608 138388 198620
rect 121236 198580 121408 198608
rect 122806 198580 138388 198608
rect 121236 198568 121242 198580
rect 97718 198500 97724 198552
rect 97776 198540 97782 198552
rect 121270 198540 121276 198552
rect 97776 198512 121276 198540
rect 97776 198500 97782 198512
rect 121270 198500 121276 198512
rect 121328 198500 121334 198552
rect 121380 198540 121408 198580
rect 138382 198568 138388 198580
rect 138440 198568 138446 198620
rect 121380 198512 132632 198540
rect 103422 198432 103428 198484
rect 103480 198472 103486 198484
rect 129734 198472 129740 198484
rect 103480 198444 129740 198472
rect 103480 198432 103486 198444
rect 129734 198432 129740 198444
rect 129792 198432 129798 198484
rect 102042 198364 102048 198416
rect 102100 198404 102106 198416
rect 126514 198404 126520 198416
rect 102100 198376 126520 198404
rect 102100 198364 102106 198376
rect 126514 198364 126520 198376
rect 126572 198364 126578 198416
rect 132604 198404 132632 198512
rect 143074 198500 143080 198552
rect 143132 198540 143138 198552
rect 146018 198540 146024 198552
rect 143132 198512 146024 198540
rect 143132 198500 143138 198512
rect 146018 198500 146024 198512
rect 146076 198500 146082 198552
rect 146588 198540 146616 198784
rect 150406 198784 164924 198812
rect 150406 198744 150434 198784
rect 173434 198772 173440 198824
rect 173492 198812 173498 198824
rect 173618 198812 173624 198824
rect 173492 198784 173624 198812
rect 173492 198772 173498 198784
rect 173618 198772 173624 198784
rect 173676 198772 173682 198824
rect 173866 198812 173894 198852
rect 174630 198840 174636 198892
rect 174688 198880 174694 198892
rect 177758 198880 177764 198892
rect 174688 198852 177764 198880
rect 174688 198840 174694 198852
rect 177758 198840 177764 198852
rect 177816 198840 177822 198892
rect 182146 198880 182174 198920
rect 185394 198880 185400 198892
rect 182146 198852 185400 198880
rect 185394 198840 185400 198852
rect 185452 198840 185458 198892
rect 178954 198812 178960 198824
rect 173866 198784 178960 198812
rect 178954 198772 178960 198784
rect 179012 198812 179018 198824
rect 179506 198812 179512 198824
rect 179012 198784 179512 198812
rect 179012 198772 179018 198784
rect 179506 198772 179512 198784
rect 179564 198772 179570 198824
rect 149026 198716 150434 198744
rect 149026 198540 149054 198716
rect 151630 198704 151636 198756
rect 151688 198744 151694 198756
rect 155218 198744 155224 198756
rect 151688 198716 155224 198744
rect 151688 198704 151694 198716
rect 155218 198704 155224 198716
rect 155276 198704 155282 198756
rect 165430 198744 165436 198756
rect 159284 198716 165436 198744
rect 150250 198636 150256 198688
rect 150308 198676 150314 198688
rect 154850 198676 154856 198688
rect 150308 198648 154856 198676
rect 150308 198636 150314 198648
rect 154850 198636 154856 198648
rect 154908 198636 154914 198688
rect 150710 198568 150716 198620
rect 150768 198608 150774 198620
rect 159284 198608 159312 198716
rect 165430 198704 165436 198716
rect 165488 198704 165494 198756
rect 167638 198704 167644 198756
rect 167696 198744 167702 198756
rect 168374 198744 168380 198756
rect 167696 198716 168380 198744
rect 167696 198704 167702 198716
rect 168374 198704 168380 198716
rect 168432 198704 168438 198756
rect 184842 198744 184848 198756
rect 169726 198716 184848 198744
rect 165614 198636 165620 198688
rect 165672 198676 165678 198688
rect 169726 198676 169754 198716
rect 184842 198704 184848 198716
rect 184900 198744 184906 198756
rect 189902 198744 189908 198756
rect 184900 198716 189908 198744
rect 184900 198704 184906 198716
rect 189902 198704 189908 198716
rect 189960 198704 189966 198756
rect 165672 198648 169754 198676
rect 165672 198636 165678 198648
rect 172974 198636 172980 198688
rect 173032 198676 173038 198688
rect 174078 198676 174084 198688
rect 173032 198648 174084 198676
rect 173032 198636 173038 198648
rect 174078 198636 174084 198648
rect 174136 198636 174142 198688
rect 182266 198636 182272 198688
rect 182324 198676 182330 198688
rect 200390 198676 200396 198688
rect 182324 198648 200396 198676
rect 182324 198636 182330 198648
rect 200390 198636 200396 198648
rect 200448 198676 200454 198688
rect 201402 198676 201408 198688
rect 200448 198648 201408 198676
rect 200448 198636 200454 198648
rect 201402 198636 201408 198648
rect 201460 198636 201466 198688
rect 150768 198580 159312 198608
rect 150768 198568 150774 198580
rect 163590 198568 163596 198620
rect 163648 198608 163654 198620
rect 169846 198608 169852 198620
rect 163648 198580 169852 198608
rect 163648 198568 163654 198580
rect 169846 198568 169852 198580
rect 169904 198568 169910 198620
rect 175642 198568 175648 198620
rect 175700 198608 175706 198620
rect 195974 198608 195980 198620
rect 175700 198580 195980 198608
rect 175700 198568 175706 198580
rect 195974 198568 195980 198580
rect 196032 198568 196038 198620
rect 146588 198512 149054 198540
rect 159726 198500 159732 198552
rect 159784 198540 159790 198552
rect 169202 198540 169208 198552
rect 159784 198512 169208 198540
rect 159784 198500 159790 198512
rect 169202 198500 169208 198512
rect 169260 198500 169266 198552
rect 171502 198500 171508 198552
rect 171560 198540 171566 198552
rect 173066 198540 173072 198552
rect 171560 198512 173072 198540
rect 171560 198500 171566 198512
rect 173066 198500 173072 198512
rect 173124 198500 173130 198552
rect 177022 198500 177028 198552
rect 177080 198540 177086 198552
rect 194502 198540 194508 198552
rect 177080 198512 194508 198540
rect 177080 198500 177086 198512
rect 194502 198500 194508 198512
rect 194560 198500 194566 198552
rect 134610 198432 134616 198484
rect 134668 198472 134674 198484
rect 140866 198472 140872 198484
rect 134668 198444 140872 198472
rect 134668 198432 134674 198444
rect 140866 198432 140872 198444
rect 140924 198432 140930 198484
rect 142430 198432 142436 198484
rect 142488 198472 142494 198484
rect 161106 198472 161112 198484
rect 142488 198444 161112 198472
rect 142488 198432 142494 198444
rect 161106 198432 161112 198444
rect 161164 198432 161170 198484
rect 161934 198432 161940 198484
rect 161992 198472 161998 198484
rect 162854 198472 162860 198484
rect 161992 198444 162860 198472
rect 161992 198432 161998 198444
rect 162854 198432 162860 198444
rect 162912 198432 162918 198484
rect 166258 198432 166264 198484
rect 166316 198472 166322 198484
rect 183554 198472 183560 198484
rect 166316 198444 183560 198472
rect 166316 198432 166322 198444
rect 183554 198432 183560 198444
rect 183612 198432 183618 198484
rect 136818 198404 136824 198416
rect 132604 198376 136824 198404
rect 136818 198364 136824 198376
rect 136876 198364 136882 198416
rect 141510 198364 141516 198416
rect 141568 198404 141574 198416
rect 147950 198404 147956 198416
rect 141568 198376 147956 198404
rect 141568 198364 141574 198376
rect 147950 198364 147956 198376
rect 148008 198364 148014 198416
rect 155862 198364 155868 198416
rect 155920 198404 155926 198416
rect 165430 198404 165436 198416
rect 155920 198376 165436 198404
rect 155920 198364 155926 198376
rect 165430 198364 165436 198376
rect 165488 198364 165494 198416
rect 165890 198364 165896 198416
rect 165948 198404 165954 198416
rect 169202 198404 169208 198416
rect 165948 198376 169208 198404
rect 165948 198364 165954 198376
rect 169202 198364 169208 198376
rect 169260 198364 169266 198416
rect 170582 198364 170588 198416
rect 170640 198404 170646 198416
rect 177666 198404 177672 198416
rect 170640 198376 177672 198404
rect 170640 198364 170646 198376
rect 177666 198364 177672 198376
rect 177724 198364 177730 198416
rect 100662 198296 100668 198348
rect 100720 198336 100726 198348
rect 133690 198336 133696 198348
rect 100720 198308 133696 198336
rect 100720 198296 100726 198308
rect 133690 198296 133696 198308
rect 133748 198296 133754 198348
rect 144086 198296 144092 198348
rect 144144 198336 144150 198348
rect 145098 198336 145104 198348
rect 144144 198308 145104 198336
rect 144144 198296 144150 198308
rect 145098 198296 145104 198308
rect 145156 198296 145162 198348
rect 156874 198296 156880 198348
rect 156932 198336 156938 198348
rect 165706 198336 165712 198348
rect 156932 198308 165712 198336
rect 156932 198296 156938 198308
rect 165706 198296 165712 198308
rect 165764 198296 165770 198348
rect 168466 198296 168472 198348
rect 168524 198336 168530 198348
rect 189258 198336 189264 198348
rect 168524 198308 189264 198336
rect 168524 198296 168530 198308
rect 189258 198296 189264 198308
rect 189316 198296 189322 198348
rect 101950 198228 101956 198280
rect 102008 198268 102014 198280
rect 134426 198268 134432 198280
rect 102008 198240 134432 198268
rect 102008 198228 102014 198240
rect 134426 198228 134432 198240
rect 134484 198228 134490 198280
rect 143552 198240 143856 198268
rect 100386 198160 100392 198212
rect 100444 198200 100450 198212
rect 126146 198200 126152 198212
rect 100444 198172 126152 198200
rect 100444 198160 100450 198172
rect 126146 198160 126152 198172
rect 126204 198160 126210 198212
rect 143552 198200 143580 198240
rect 137986 198172 143580 198200
rect 143828 198200 143856 198240
rect 148042 198228 148048 198280
rect 148100 198268 148106 198280
rect 148410 198268 148416 198280
rect 148100 198240 148416 198268
rect 148100 198228 148106 198240
rect 148410 198228 148416 198240
rect 148468 198268 148474 198280
rect 169018 198268 169024 198280
rect 148468 198240 169024 198268
rect 148468 198228 148474 198240
rect 169018 198228 169024 198240
rect 169076 198228 169082 198280
rect 169202 198228 169208 198280
rect 169260 198268 169266 198280
rect 189166 198268 189172 198280
rect 169260 198240 189172 198268
rect 169260 198228 169266 198240
rect 189166 198228 189172 198240
rect 189224 198228 189230 198280
rect 164234 198200 164240 198212
rect 143828 198172 145696 198200
rect 106182 198092 106188 198144
rect 106240 198132 106246 198144
rect 106240 198104 133184 198132
rect 106240 198092 106246 198104
rect 100570 198024 100576 198076
rect 100628 198064 100634 198076
rect 100628 198036 131896 198064
rect 100628 198024 100634 198036
rect 61378 197956 61384 198008
rect 61436 197996 61442 198008
rect 99282 197996 99288 198008
rect 61436 197968 99288 197996
rect 61436 197956 61442 197968
rect 99282 197956 99288 197968
rect 99340 197996 99346 198008
rect 127158 197996 127164 198008
rect 99340 197968 127164 197996
rect 99340 197956 99346 197968
rect 127158 197956 127164 197968
rect 127216 197956 127222 198008
rect 122190 197888 122196 197940
rect 122248 197928 122254 197940
rect 131758 197928 131764 197940
rect 122248 197900 131764 197928
rect 122248 197888 122254 197900
rect 131758 197888 131764 197900
rect 131816 197888 131822 197940
rect 131868 197928 131896 198036
rect 133156 197996 133184 198104
rect 135990 198024 135996 198076
rect 136048 198064 136054 198076
rect 137986 198064 138014 198172
rect 142246 198092 142252 198144
rect 142304 198132 142310 198144
rect 143442 198132 143448 198144
rect 142304 198104 143448 198132
rect 142304 198092 142310 198104
rect 143442 198092 143448 198104
rect 143500 198092 143506 198144
rect 136048 198036 138014 198064
rect 145668 198064 145696 198172
rect 164206 198160 164240 198200
rect 164292 198160 164298 198212
rect 171778 198160 171784 198212
rect 171836 198200 171842 198212
rect 172974 198200 172980 198212
rect 171836 198172 172980 198200
rect 171836 198160 171842 198172
rect 172974 198160 172980 198172
rect 173032 198160 173038 198212
rect 178402 198160 178408 198212
rect 178460 198200 178466 198212
rect 208394 198200 208400 198212
rect 178460 198172 208400 198200
rect 178460 198160 178466 198172
rect 208394 198160 208400 198172
rect 208452 198160 208458 198212
rect 152918 198092 152924 198144
rect 152976 198132 152982 198144
rect 154666 198132 154672 198144
rect 152976 198104 154672 198132
rect 152976 198092 152982 198104
rect 154666 198092 154672 198104
rect 154724 198092 154730 198144
rect 155954 198092 155960 198144
rect 156012 198132 156018 198144
rect 164206 198132 164234 198160
rect 169294 198132 169300 198144
rect 156012 198104 164234 198132
rect 167196 198104 169300 198132
rect 156012 198092 156018 198104
rect 162762 198064 162768 198076
rect 145668 198036 162768 198064
rect 136048 198024 136054 198036
rect 162762 198024 162768 198036
rect 162820 198024 162826 198076
rect 165430 198024 165436 198076
rect 165488 198064 165494 198076
rect 167196 198064 167224 198104
rect 169294 198092 169300 198104
rect 169352 198092 169358 198144
rect 172238 198092 172244 198144
rect 172296 198132 172302 198144
rect 173894 198132 173900 198144
rect 172296 198104 173900 198132
rect 172296 198092 172302 198104
rect 173894 198092 173900 198104
rect 173952 198092 173958 198144
rect 182174 198092 182180 198144
rect 182232 198132 182238 198144
rect 219526 198132 219532 198144
rect 182232 198104 219532 198132
rect 182232 198092 182238 198104
rect 219526 198092 219532 198104
rect 219584 198132 219590 198144
rect 220722 198132 220728 198144
rect 219584 198104 220728 198132
rect 219584 198092 219590 198104
rect 220722 198092 220728 198104
rect 220780 198092 220786 198144
rect 165488 198036 167224 198064
rect 165488 198024 165494 198036
rect 169386 198024 169392 198076
rect 169444 198064 169450 198076
rect 219434 198064 219440 198076
rect 169444 198036 219440 198064
rect 169444 198024 169450 198036
rect 219434 198024 219440 198036
rect 219492 198024 219498 198076
rect 138014 197996 138020 198008
rect 133156 197968 138020 197996
rect 138014 197956 138020 197968
rect 138072 197956 138078 198008
rect 143442 197956 143448 198008
rect 143500 197996 143506 198008
rect 146938 197996 146944 198008
rect 143500 197968 146944 197996
rect 143500 197956 143506 197968
rect 146938 197956 146944 197968
rect 146996 197956 147002 198008
rect 561306 197996 561312 198008
rect 158180 197968 561312 197996
rect 133966 197928 133972 197940
rect 131868 197900 133972 197928
rect 133966 197888 133972 197900
rect 134024 197888 134030 197940
rect 139578 197888 139584 197940
rect 139636 197928 139642 197940
rect 144178 197928 144184 197940
rect 139636 197900 144184 197928
rect 139636 197888 139642 197900
rect 144178 197888 144184 197900
rect 144236 197928 144242 197940
rect 158180 197928 158208 197968
rect 561306 197956 561312 197968
rect 561364 197956 561370 198008
rect 144236 197900 158208 197928
rect 144236 197888 144242 197900
rect 162946 197888 162952 197940
rect 163004 197928 163010 197940
rect 177482 197928 177488 197940
rect 163004 197900 177488 197928
rect 163004 197888 163010 197900
rect 177482 197888 177488 197900
rect 177540 197888 177546 197940
rect 138750 197820 138756 197872
rect 138808 197860 138814 197872
rect 145926 197860 145932 197872
rect 138808 197832 145932 197860
rect 138808 197820 138814 197832
rect 145926 197820 145932 197832
rect 145984 197820 145990 197872
rect 152090 197820 152096 197872
rect 152148 197860 152154 197872
rect 154758 197860 154764 197872
rect 152148 197832 154764 197860
rect 152148 197820 152154 197832
rect 154758 197820 154764 197832
rect 154816 197820 154822 197872
rect 127802 197752 127808 197804
rect 127860 197792 127866 197804
rect 138198 197792 138204 197804
rect 127860 197764 138204 197792
rect 127860 197752 127866 197764
rect 138198 197752 138204 197764
rect 138256 197752 138262 197804
rect 145558 197752 145564 197804
rect 145616 197792 145622 197804
rect 148226 197792 148232 197804
rect 145616 197764 148232 197792
rect 145616 197752 145622 197764
rect 148226 197752 148232 197764
rect 148284 197752 148290 197804
rect 149054 197752 149060 197804
rect 149112 197792 149118 197804
rect 149112 197764 156092 197792
rect 149112 197752 149118 197764
rect 113174 197684 113180 197736
rect 113232 197724 113238 197736
rect 131022 197724 131028 197736
rect 113232 197696 131028 197724
rect 113232 197684 113238 197696
rect 131022 197684 131028 197696
rect 131080 197684 131086 197736
rect 141418 197684 141424 197736
rect 141476 197724 141482 197736
rect 149072 197724 149100 197752
rect 141476 197696 149100 197724
rect 141476 197684 141482 197696
rect 133138 197616 133144 197668
rect 133196 197656 133202 197668
rect 142614 197656 142620 197668
rect 133196 197628 142620 197656
rect 133196 197616 133202 197628
rect 142614 197616 142620 197628
rect 142672 197616 142678 197668
rect 148042 197616 148048 197668
rect 148100 197656 148106 197668
rect 150802 197656 150808 197668
rect 148100 197628 150808 197656
rect 148100 197616 148106 197628
rect 150802 197616 150808 197628
rect 150860 197616 150866 197668
rect 133966 197548 133972 197600
rect 134024 197588 134030 197600
rect 144454 197588 144460 197600
rect 134024 197560 144460 197588
rect 134024 197548 134030 197560
rect 144454 197548 144460 197560
rect 144512 197548 144518 197600
rect 156064 197588 156092 197764
rect 160278 197752 160284 197804
rect 160336 197792 160342 197804
rect 169386 197792 169392 197804
rect 160336 197764 169392 197792
rect 160336 197752 160342 197764
rect 169386 197752 169392 197764
rect 169444 197752 169450 197804
rect 177574 197752 177580 197804
rect 177632 197792 177638 197804
rect 178218 197792 178224 197804
rect 177632 197764 178224 197792
rect 177632 197752 177638 197764
rect 178218 197752 178224 197764
rect 178276 197752 178282 197804
rect 157150 197684 157156 197736
rect 157208 197724 157214 197736
rect 164234 197724 164240 197736
rect 157208 197696 164240 197724
rect 157208 197684 157214 197696
rect 164234 197684 164240 197696
rect 164292 197684 164298 197736
rect 172514 197684 172520 197736
rect 172572 197724 172578 197736
rect 172882 197724 172888 197736
rect 172572 197696 172888 197724
rect 172572 197684 172578 197696
rect 172882 197684 172888 197696
rect 172940 197684 172946 197736
rect 161842 197616 161848 197668
rect 161900 197656 161906 197668
rect 170582 197656 170588 197668
rect 161900 197628 170588 197656
rect 161900 197616 161906 197628
rect 170582 197616 170588 197628
rect 170640 197616 170646 197668
rect 171410 197616 171416 197668
rect 171468 197656 171474 197668
rect 177574 197656 177580 197668
rect 171468 197628 177580 197656
rect 171468 197616 171474 197628
rect 177574 197616 177580 197628
rect 177632 197616 177638 197668
rect 170766 197588 170772 197600
rect 156064 197560 170772 197588
rect 170766 197548 170772 197560
rect 170824 197548 170830 197600
rect 138014 197480 138020 197532
rect 138072 197520 138078 197532
rect 138750 197520 138756 197532
rect 138072 197492 138756 197520
rect 138072 197480 138078 197492
rect 138750 197480 138756 197492
rect 138808 197480 138814 197532
rect 140038 197480 140044 197532
rect 140096 197520 140102 197532
rect 147858 197520 147864 197532
rect 140096 197492 147864 197520
rect 140096 197480 140102 197492
rect 147858 197480 147864 197492
rect 147916 197480 147922 197532
rect 151630 197480 151636 197532
rect 151688 197520 151694 197532
rect 153930 197520 153936 197532
rect 151688 197492 153936 197520
rect 151688 197480 151694 197492
rect 153930 197480 153936 197492
rect 153988 197480 153994 197532
rect 154942 197480 154948 197532
rect 155000 197520 155006 197532
rect 155402 197520 155408 197532
rect 155000 197492 155408 197520
rect 155000 197480 155006 197492
rect 155402 197480 155408 197492
rect 155460 197480 155466 197532
rect 160830 197480 160836 197532
rect 160888 197520 160894 197532
rect 165614 197520 165620 197532
rect 160888 197492 165620 197520
rect 160888 197480 160894 197492
rect 165614 197480 165620 197492
rect 165672 197480 165678 197532
rect 146754 197412 146760 197464
rect 146812 197452 146818 197464
rect 147306 197452 147312 197464
rect 146812 197424 147312 197452
rect 146812 197412 146818 197424
rect 147306 197412 147312 197424
rect 147364 197412 147370 197464
rect 149054 197412 149060 197464
rect 149112 197452 149118 197464
rect 150342 197452 150348 197464
rect 149112 197424 150348 197452
rect 149112 197412 149118 197424
rect 150342 197412 150348 197424
rect 150400 197412 150406 197464
rect 164970 197412 164976 197464
rect 165028 197452 165034 197464
rect 168006 197452 168012 197464
rect 165028 197424 168012 197452
rect 165028 197412 165034 197424
rect 168006 197412 168012 197424
rect 168064 197412 168070 197464
rect 139486 197344 139492 197396
rect 139544 197384 139550 197396
rect 143810 197384 143816 197396
rect 139544 197356 143816 197384
rect 139544 197344 139550 197356
rect 143810 197344 143816 197356
rect 143868 197344 143874 197396
rect 146662 197344 146668 197396
rect 146720 197384 146726 197396
rect 147122 197384 147128 197396
rect 146720 197356 147128 197384
rect 146720 197344 146726 197356
rect 147122 197344 147128 197356
rect 147180 197344 147186 197396
rect 147950 197344 147956 197396
rect 148008 197384 148014 197396
rect 150710 197384 150716 197396
rect 148008 197356 150716 197384
rect 148008 197344 148014 197356
rect 150710 197344 150716 197356
rect 150768 197344 150774 197396
rect 168650 197344 168656 197396
rect 168708 197384 168714 197396
rect 171502 197384 171508 197396
rect 168708 197356 171508 197384
rect 168708 197344 168714 197356
rect 171502 197344 171508 197356
rect 171560 197344 171566 197396
rect 172698 197344 172704 197396
rect 172756 197384 172762 197396
rect 172756 197356 176654 197384
rect 172756 197344 172762 197356
rect 108390 197276 108396 197328
rect 108448 197316 108454 197328
rect 170858 197316 170864 197328
rect 108448 197288 170864 197316
rect 108448 197276 108454 197288
rect 170858 197276 170864 197288
rect 170916 197276 170922 197328
rect 176626 197316 176654 197356
rect 220722 197344 220728 197396
rect 220780 197384 220786 197396
rect 580166 197384 580172 197396
rect 220780 197356 580172 197384
rect 220780 197344 220786 197356
rect 580166 197344 580172 197356
rect 580224 197344 580230 197396
rect 192294 197316 192300 197328
rect 176626 197288 192300 197316
rect 192294 197276 192300 197288
rect 192352 197316 192358 197328
rect 193122 197316 193128 197328
rect 192352 197288 193128 197316
rect 192352 197276 192358 197288
rect 193122 197276 193128 197288
rect 193180 197276 193186 197328
rect 97350 197208 97356 197260
rect 97408 197248 97414 197260
rect 161382 197248 161388 197260
rect 97408 197220 161388 197248
rect 97408 197208 97414 197220
rect 161382 197208 161388 197220
rect 161440 197248 161446 197260
rect 164050 197248 164056 197260
rect 161440 197220 164056 197248
rect 161440 197208 161446 197220
rect 164050 197208 164056 197220
rect 164108 197208 164114 197260
rect 170766 197248 170772 197260
rect 164206 197220 170772 197248
rect 111150 197140 111156 197192
rect 111208 197180 111214 197192
rect 164206 197180 164234 197220
rect 170766 197208 170772 197220
rect 170824 197248 170830 197260
rect 171962 197248 171968 197260
rect 170824 197220 171968 197248
rect 170824 197208 170830 197220
rect 171962 197208 171968 197220
rect 172020 197208 172026 197260
rect 172330 197208 172336 197260
rect 172388 197248 172394 197260
rect 173342 197248 173348 197260
rect 172388 197220 173348 197248
rect 172388 197208 172394 197220
rect 173342 197208 173348 197220
rect 173400 197208 173406 197260
rect 173894 197208 173900 197260
rect 173952 197248 173958 197260
rect 189626 197248 189632 197260
rect 173952 197220 189632 197248
rect 173952 197208 173958 197220
rect 189626 197208 189632 197220
rect 189684 197248 189690 197260
rect 209866 197248 209872 197260
rect 189684 197220 209872 197248
rect 189684 197208 189690 197220
rect 209866 197208 209872 197220
rect 209924 197208 209930 197260
rect 111208 197152 164234 197180
rect 111208 197140 111214 197152
rect 169754 197140 169760 197192
rect 169812 197180 169818 197192
rect 171410 197180 171416 197192
rect 169812 197152 171416 197180
rect 169812 197140 169818 197152
rect 171410 197140 171416 197152
rect 171468 197140 171474 197192
rect 171594 197140 171600 197192
rect 171652 197180 171658 197192
rect 192570 197180 192576 197192
rect 171652 197152 192576 197180
rect 171652 197140 171658 197152
rect 192570 197140 192576 197152
rect 192628 197140 192634 197192
rect 112438 197072 112444 197124
rect 112496 197112 112502 197124
rect 112496 197084 138014 197112
rect 112496 197072 112502 197084
rect 104250 197004 104256 197056
rect 104308 197044 104314 197056
rect 107286 197044 107292 197056
rect 104308 197016 107292 197044
rect 104308 197004 104314 197016
rect 107286 197004 107292 197016
rect 107344 197044 107350 197056
rect 132402 197044 132408 197056
rect 107344 197016 132408 197044
rect 107344 197004 107350 197016
rect 132402 197004 132408 197016
rect 132460 197004 132466 197056
rect 135898 197004 135904 197056
rect 135956 197044 135962 197056
rect 136358 197044 136364 197056
rect 135956 197016 136364 197044
rect 135956 197004 135962 197016
rect 136358 197004 136364 197016
rect 136416 197004 136422 197056
rect 136450 197004 136456 197056
rect 136508 197044 136514 197056
rect 136634 197044 136640 197056
rect 136508 197016 136640 197044
rect 136508 197004 136514 197016
rect 136634 197004 136640 197016
rect 136692 197004 136698 197056
rect 137986 197044 138014 197084
rect 146662 197072 146668 197124
rect 146720 197112 146726 197124
rect 148134 197112 148140 197124
rect 146720 197084 148140 197112
rect 146720 197072 146726 197084
rect 148134 197072 148140 197084
rect 148192 197072 148198 197124
rect 149238 197072 149244 197124
rect 149296 197112 149302 197124
rect 149698 197112 149704 197124
rect 149296 197084 149704 197112
rect 149296 197072 149302 197084
rect 149698 197072 149704 197084
rect 149756 197072 149762 197124
rect 149790 197072 149796 197124
rect 149848 197112 149854 197124
rect 150342 197112 150348 197124
rect 149848 197084 150348 197112
rect 149848 197072 149854 197084
rect 150342 197072 150348 197084
rect 150400 197072 150406 197124
rect 161474 197072 161480 197124
rect 161532 197112 161538 197124
rect 191926 197112 191932 197124
rect 161532 197084 191932 197112
rect 161532 197072 161538 197084
rect 191926 197072 191932 197084
rect 191984 197072 191990 197124
rect 193122 197072 193128 197124
rect 193180 197112 193186 197124
rect 209958 197112 209964 197124
rect 193180 197084 209964 197112
rect 193180 197072 193186 197084
rect 209958 197072 209964 197084
rect 210016 197072 210022 197124
rect 137986 197016 154574 197044
rect 118326 196936 118332 196988
rect 118384 196976 118390 196988
rect 149514 196976 149520 196988
rect 118384 196948 149520 196976
rect 118384 196936 118390 196948
rect 149514 196936 149520 196948
rect 149572 196936 149578 196988
rect 153102 196936 153108 196988
rect 153160 196976 153166 196988
rect 153838 196976 153844 196988
rect 153160 196948 153844 196976
rect 153160 196936 153166 196948
rect 153838 196936 153844 196948
rect 153896 196936 153902 196988
rect 154546 196976 154574 197016
rect 158530 197004 158536 197056
rect 158588 197044 158594 197056
rect 159634 197044 159640 197056
rect 158588 197016 159640 197044
rect 158588 197004 158594 197016
rect 159634 197004 159640 197016
rect 159692 197004 159698 197056
rect 166074 197004 166080 197056
rect 166132 197044 166138 197056
rect 200206 197044 200212 197056
rect 166132 197016 200212 197044
rect 166132 197004 166138 197016
rect 200206 197004 200212 197016
rect 200264 197004 200270 197056
rect 156414 196976 156420 196988
rect 154546 196948 156420 196976
rect 156414 196936 156420 196948
rect 156472 196976 156478 196988
rect 171870 196976 171876 196988
rect 156472 196948 171876 196976
rect 156472 196936 156478 196948
rect 171870 196936 171876 196948
rect 171928 196936 171934 196988
rect 171962 196936 171968 196988
rect 172020 196976 172026 196988
rect 208486 196976 208492 196988
rect 172020 196948 208492 196976
rect 172020 196936 172026 196948
rect 208486 196936 208492 196948
rect 208544 196936 208550 196988
rect 104802 196868 104808 196920
rect 104860 196908 104866 196920
rect 138566 196908 138572 196920
rect 104860 196880 138572 196908
rect 104860 196868 104866 196880
rect 138566 196868 138572 196880
rect 138624 196868 138630 196920
rect 144822 196868 144828 196920
rect 144880 196908 144886 196920
rect 147030 196908 147036 196920
rect 144880 196880 147036 196908
rect 144880 196868 144886 196880
rect 147030 196868 147036 196880
rect 147088 196868 147094 196920
rect 148318 196868 148324 196920
rect 148376 196908 148382 196920
rect 148502 196908 148508 196920
rect 148376 196880 148508 196908
rect 148376 196868 148382 196880
rect 148502 196868 148508 196880
rect 148560 196868 148566 196920
rect 157242 196868 157248 196920
rect 157300 196908 157306 196920
rect 157518 196908 157524 196920
rect 157300 196880 157524 196908
rect 157300 196868 157306 196880
rect 157518 196868 157524 196880
rect 157576 196868 157582 196920
rect 170306 196908 170312 196920
rect 159284 196880 170312 196908
rect 158162 196840 158168 196852
rect 122806 196812 158168 196840
rect 117958 196732 117964 196784
rect 118016 196772 118022 196784
rect 122806 196772 122834 196812
rect 158162 196800 158168 196812
rect 158220 196800 158226 196852
rect 158254 196800 158260 196852
rect 158312 196840 158318 196852
rect 159284 196840 159312 196880
rect 170306 196868 170312 196880
rect 170364 196868 170370 196920
rect 170858 196868 170864 196920
rect 170916 196908 170922 196920
rect 174078 196908 174084 196920
rect 170916 196880 174084 196908
rect 170916 196868 170922 196880
rect 174078 196868 174084 196880
rect 174136 196908 174142 196920
rect 212718 196908 212724 196920
rect 174136 196880 212724 196908
rect 174136 196868 174142 196880
rect 212718 196868 212724 196880
rect 212776 196868 212782 196920
rect 158312 196812 159312 196840
rect 158312 196800 158318 196812
rect 159358 196800 159364 196852
rect 159416 196840 159422 196852
rect 163498 196840 163504 196852
rect 159416 196812 163504 196840
rect 159416 196800 159422 196812
rect 163498 196800 163504 196812
rect 163556 196800 163562 196852
rect 167914 196800 167920 196852
rect 167972 196840 167978 196852
rect 169202 196840 169208 196852
rect 167972 196812 169208 196840
rect 167972 196800 167978 196812
rect 169202 196800 169208 196812
rect 169260 196800 169266 196852
rect 170766 196800 170772 196852
rect 170824 196840 170830 196852
rect 173342 196840 173348 196852
rect 170824 196812 173348 196840
rect 170824 196800 170830 196812
rect 173342 196800 173348 196812
rect 173400 196840 173406 196852
rect 212626 196840 212632 196852
rect 173400 196812 212632 196840
rect 173400 196800 173406 196812
rect 212626 196800 212632 196812
rect 212684 196800 212690 196852
rect 118016 196744 122834 196772
rect 118016 196732 118022 196744
rect 138750 196732 138756 196784
rect 138808 196772 138814 196784
rect 141050 196772 141056 196784
rect 138808 196744 141056 196772
rect 138808 196732 138814 196744
rect 141050 196732 141056 196744
rect 141108 196732 141114 196784
rect 143534 196732 143540 196784
rect 143592 196772 143598 196784
rect 144454 196772 144460 196784
rect 143592 196744 144460 196772
rect 143592 196732 143598 196744
rect 144454 196732 144460 196744
rect 144512 196732 144518 196784
rect 146386 196732 146392 196784
rect 146444 196772 146450 196784
rect 146846 196772 146852 196784
rect 146444 196744 146852 196772
rect 146444 196732 146450 196744
rect 146846 196732 146852 196744
rect 146904 196732 146910 196784
rect 148134 196732 148140 196784
rect 148192 196772 148198 196784
rect 148778 196772 148784 196784
rect 148192 196744 148784 196772
rect 148192 196732 148198 196744
rect 148778 196732 148784 196744
rect 148836 196732 148842 196784
rect 154666 196732 154672 196784
rect 154724 196772 154730 196784
rect 155586 196772 155592 196784
rect 154724 196744 155592 196772
rect 154724 196732 154730 196744
rect 155586 196732 155592 196744
rect 155644 196732 155650 196784
rect 155678 196732 155684 196784
rect 155736 196772 155742 196784
rect 155862 196772 155868 196784
rect 155736 196744 155868 196772
rect 155736 196732 155742 196744
rect 155862 196732 155868 196744
rect 155920 196732 155926 196784
rect 156138 196732 156144 196784
rect 156196 196772 156202 196784
rect 156782 196772 156788 196784
rect 156196 196744 156788 196772
rect 156196 196732 156202 196744
rect 156782 196732 156788 196744
rect 156840 196732 156846 196784
rect 157518 196732 157524 196784
rect 157576 196772 157582 196784
rect 158346 196772 158352 196784
rect 157576 196744 158352 196772
rect 157576 196732 157582 196744
rect 158346 196732 158352 196744
rect 158404 196732 158410 196784
rect 158990 196732 158996 196784
rect 159048 196772 159054 196784
rect 160002 196772 160008 196784
rect 159048 196744 160008 196772
rect 159048 196732 159054 196744
rect 160002 196732 160008 196744
rect 160060 196732 160066 196784
rect 163130 196732 163136 196784
rect 163188 196772 163194 196784
rect 214650 196772 214656 196784
rect 163188 196744 214656 196772
rect 163188 196732 163194 196744
rect 214650 196732 214656 196744
rect 214708 196732 214714 196784
rect 96522 196664 96528 196716
rect 96580 196704 96586 196716
rect 124398 196704 124404 196716
rect 96580 196676 124404 196704
rect 96580 196664 96586 196676
rect 124398 196664 124404 196676
rect 124456 196664 124462 196716
rect 136358 196664 136364 196716
rect 136416 196704 136422 196716
rect 136634 196704 136640 196716
rect 136416 196676 136640 196704
rect 136416 196664 136422 196676
rect 136634 196664 136640 196676
rect 136692 196664 136698 196716
rect 139578 196664 139584 196716
rect 139636 196704 139642 196716
rect 140682 196704 140688 196716
rect 139636 196676 140688 196704
rect 139636 196664 139642 196676
rect 140682 196664 140688 196676
rect 140740 196664 140746 196716
rect 141970 196664 141976 196716
rect 142028 196704 142034 196716
rect 143166 196704 143172 196716
rect 142028 196676 143172 196704
rect 142028 196664 142034 196676
rect 143166 196664 143172 196676
rect 143224 196664 143230 196716
rect 143718 196664 143724 196716
rect 143776 196704 143782 196716
rect 144270 196704 144276 196716
rect 143776 196676 144276 196704
rect 143776 196664 143782 196676
rect 144270 196664 144276 196676
rect 144328 196664 144334 196716
rect 146754 196664 146760 196716
rect 146812 196704 146818 196716
rect 147582 196704 147588 196716
rect 146812 196676 147588 196704
rect 146812 196664 146818 196676
rect 147582 196664 147588 196676
rect 147640 196664 147646 196716
rect 147674 196664 147680 196716
rect 147732 196704 147738 196716
rect 148870 196704 148876 196716
rect 147732 196676 148876 196704
rect 147732 196664 147738 196676
rect 148870 196664 148876 196676
rect 148928 196664 148934 196716
rect 149514 196664 149520 196716
rect 149572 196704 149578 196716
rect 150066 196704 150072 196716
rect 149572 196676 150072 196704
rect 149572 196664 149578 196676
rect 150066 196664 150072 196676
rect 150124 196664 150130 196716
rect 150526 196664 150532 196716
rect 150584 196704 150590 196716
rect 151446 196704 151452 196716
rect 150584 196676 151452 196704
rect 150584 196664 150590 196676
rect 151446 196664 151452 196676
rect 151504 196664 151510 196716
rect 152826 196664 152832 196716
rect 152884 196704 152890 196716
rect 215294 196704 215300 196716
rect 152884 196676 215300 196704
rect 152884 196664 152890 196676
rect 215294 196664 215300 196676
rect 215352 196664 215358 196716
rect 3142 196596 3148 196648
rect 3200 196636 3206 196648
rect 167270 196636 167276 196648
rect 3200 196608 167276 196636
rect 3200 196596 3206 196608
rect 167270 196596 167276 196608
rect 167328 196636 167334 196648
rect 169018 196636 169024 196648
rect 167328 196608 169024 196636
rect 167328 196596 167334 196608
rect 169018 196596 169024 196608
rect 169076 196596 169082 196648
rect 169754 196596 169760 196648
rect 169812 196636 169818 196648
rect 170030 196636 170036 196648
rect 169812 196608 170036 196636
rect 169812 196596 169818 196608
rect 170030 196596 170036 196608
rect 170088 196596 170094 196648
rect 170490 196596 170496 196648
rect 170548 196636 170554 196648
rect 173342 196636 173348 196648
rect 170548 196608 173348 196636
rect 170548 196596 170554 196608
rect 173342 196596 173348 196608
rect 173400 196596 173406 196648
rect 174078 196596 174084 196648
rect 174136 196636 174142 196648
rect 174354 196636 174360 196648
rect 174136 196608 174360 196636
rect 174136 196596 174142 196608
rect 174354 196596 174360 196608
rect 174412 196596 174418 196648
rect 185394 196596 185400 196648
rect 185452 196636 185458 196648
rect 207106 196636 207112 196648
rect 185452 196608 207112 196636
rect 185452 196596 185458 196608
rect 207106 196596 207112 196608
rect 207164 196636 207170 196648
rect 563698 196636 563704 196648
rect 207164 196608 563704 196636
rect 207164 196596 207170 196608
rect 563698 196596 563704 196608
rect 563756 196596 563762 196648
rect 121270 196528 121276 196580
rect 121328 196568 121334 196580
rect 125410 196568 125416 196580
rect 121328 196540 125416 196568
rect 121328 196528 121334 196540
rect 125410 196528 125416 196540
rect 125468 196528 125474 196580
rect 142154 196528 142160 196580
rect 142212 196568 142218 196580
rect 144730 196568 144736 196580
rect 142212 196540 144736 196568
rect 142212 196528 142218 196540
rect 144730 196528 144736 196540
rect 144788 196528 144794 196580
rect 145190 196528 145196 196580
rect 145248 196568 145254 196580
rect 145834 196568 145840 196580
rect 145248 196540 145840 196568
rect 145248 196528 145254 196540
rect 145834 196528 145840 196540
rect 145892 196528 145898 196580
rect 154850 196528 154856 196580
rect 154908 196568 154914 196580
rect 155770 196568 155776 196580
rect 154908 196540 155776 196568
rect 154908 196528 154914 196540
rect 155770 196528 155776 196540
rect 155828 196528 155834 196580
rect 159082 196528 159088 196580
rect 159140 196568 159146 196580
rect 159542 196568 159548 196580
rect 159140 196540 159548 196568
rect 159140 196528 159146 196540
rect 159542 196528 159548 196540
rect 159600 196528 159606 196580
rect 160186 196528 160192 196580
rect 160244 196568 160250 196580
rect 160370 196568 160376 196580
rect 160244 196540 160376 196568
rect 160244 196528 160250 196540
rect 160370 196528 160376 196540
rect 160428 196528 160434 196580
rect 163682 196528 163688 196580
rect 163740 196568 163746 196580
rect 164142 196568 164148 196580
rect 163740 196540 164148 196568
rect 163740 196528 163746 196540
rect 164142 196528 164148 196540
rect 164200 196528 164206 196580
rect 168466 196528 168472 196580
rect 168524 196568 168530 196580
rect 169478 196568 169484 196580
rect 168524 196540 169484 196568
rect 168524 196528 168530 196540
rect 169478 196528 169484 196540
rect 169536 196528 169542 196580
rect 170122 196528 170128 196580
rect 170180 196568 170186 196580
rect 171962 196568 171968 196580
rect 170180 196540 171968 196568
rect 170180 196528 170186 196540
rect 171962 196528 171968 196540
rect 172020 196528 172026 196580
rect 131850 196460 131856 196512
rect 131908 196500 131914 196512
rect 140774 196500 140780 196512
rect 131908 196472 140780 196500
rect 131908 196460 131914 196472
rect 140774 196460 140780 196472
rect 140832 196460 140838 196512
rect 143718 196460 143724 196512
rect 143776 196500 143782 196512
rect 144638 196500 144644 196512
rect 143776 196472 144644 196500
rect 143776 196460 143782 196472
rect 144638 196460 144644 196472
rect 144696 196460 144702 196512
rect 150710 196460 150716 196512
rect 150768 196500 150774 196512
rect 151354 196500 151360 196512
rect 150768 196472 151360 196500
rect 150768 196460 150774 196472
rect 151354 196460 151360 196472
rect 151412 196460 151418 196512
rect 155034 196460 155040 196512
rect 155092 196500 155098 196512
rect 155586 196500 155592 196512
rect 155092 196472 155592 196500
rect 155092 196460 155098 196472
rect 155586 196460 155592 196472
rect 155644 196460 155650 196512
rect 156046 196460 156052 196512
rect 156104 196500 156110 196512
rect 156874 196500 156880 196512
rect 156104 196472 156880 196500
rect 156104 196460 156110 196472
rect 156874 196460 156880 196472
rect 156932 196460 156938 196512
rect 157702 196460 157708 196512
rect 157760 196500 157766 196512
rect 160830 196500 160836 196512
rect 157760 196472 160836 196500
rect 157760 196460 157766 196472
rect 160830 196460 160836 196472
rect 160888 196460 160894 196512
rect 164050 196460 164056 196512
rect 164108 196500 164114 196512
rect 178678 196500 178684 196512
rect 164108 196472 178684 196500
rect 164108 196460 164114 196472
rect 178678 196460 178684 196472
rect 178736 196460 178742 196512
rect 116486 196392 116492 196444
rect 116544 196432 116550 196444
rect 116544 196404 138014 196432
rect 116544 196392 116550 196404
rect 137986 196364 138014 196404
rect 141602 196392 141608 196444
rect 141660 196432 141666 196444
rect 142430 196432 142436 196444
rect 141660 196404 142436 196432
rect 141660 196392 141666 196404
rect 142430 196392 142436 196404
rect 142488 196392 142494 196444
rect 144914 196392 144920 196444
rect 144972 196432 144978 196444
rect 145834 196432 145840 196444
rect 144972 196404 145840 196432
rect 144972 196392 144978 196404
rect 145834 196392 145840 196404
rect 145892 196392 145898 196444
rect 158070 196392 158076 196444
rect 158128 196432 158134 196444
rect 158530 196432 158536 196444
rect 158128 196404 158536 196432
rect 158128 196392 158134 196404
rect 158530 196392 158536 196404
rect 158588 196392 158594 196444
rect 161658 196432 161664 196444
rect 159054 196404 161664 196432
rect 159054 196364 159082 196404
rect 161658 196392 161664 196404
rect 161716 196392 161722 196444
rect 162946 196392 162952 196444
rect 163004 196432 163010 196444
rect 163958 196432 163964 196444
rect 163004 196404 163964 196432
rect 163004 196392 163010 196404
rect 163958 196392 163964 196404
rect 164016 196392 164022 196444
rect 164418 196392 164424 196444
rect 164476 196432 164482 196444
rect 164694 196432 164700 196444
rect 164476 196404 164700 196432
rect 164476 196392 164482 196404
rect 164694 196392 164700 196404
rect 164752 196392 164758 196444
rect 165982 196392 165988 196444
rect 166040 196432 166046 196444
rect 166810 196432 166816 196444
rect 166040 196404 166816 196432
rect 166040 196392 166046 196404
rect 166810 196392 166816 196404
rect 166868 196392 166874 196444
rect 168558 196392 168564 196444
rect 168616 196432 168622 196444
rect 168926 196432 168932 196444
rect 168616 196404 168932 196432
rect 168616 196392 168622 196404
rect 168926 196392 168932 196404
rect 168984 196392 168990 196444
rect 171134 196392 171140 196444
rect 171192 196432 171198 196444
rect 172054 196432 172060 196444
rect 171192 196404 172060 196432
rect 171192 196392 171198 196404
rect 172054 196392 172060 196404
rect 172112 196392 172118 196444
rect 176286 196392 176292 196444
rect 176344 196432 176350 196444
rect 178402 196432 178408 196444
rect 176344 196404 178408 196432
rect 176344 196392 176350 196404
rect 178402 196392 178408 196404
rect 178460 196392 178466 196444
rect 137986 196336 159082 196364
rect 166994 196324 167000 196376
rect 167052 196364 167058 196376
rect 172882 196364 172888 196376
rect 167052 196336 172888 196364
rect 167052 196324 167058 196336
rect 172882 196324 172888 196336
rect 172940 196324 172946 196376
rect 131942 196256 131948 196308
rect 132000 196296 132006 196308
rect 138934 196296 138940 196308
rect 132000 196268 138940 196296
rect 132000 196256 132006 196268
rect 138934 196256 138940 196268
rect 138992 196256 138998 196308
rect 140314 196256 140320 196308
rect 140372 196296 140378 196308
rect 141602 196296 141608 196308
rect 140372 196268 141608 196296
rect 140372 196256 140378 196268
rect 141602 196256 141608 196268
rect 141660 196256 141666 196308
rect 156598 196256 156604 196308
rect 156656 196296 156662 196308
rect 156966 196296 156972 196308
rect 156656 196268 156972 196296
rect 156656 196256 156662 196268
rect 156966 196256 156972 196268
rect 157024 196256 157030 196308
rect 159450 196256 159456 196308
rect 159508 196296 159514 196308
rect 173158 196296 173164 196308
rect 159508 196268 173164 196296
rect 159508 196256 159514 196268
rect 173158 196256 173164 196268
rect 173216 196256 173222 196308
rect 158162 196188 158168 196240
rect 158220 196228 158226 196240
rect 159726 196228 159732 196240
rect 158220 196200 159732 196228
rect 158220 196188 158226 196200
rect 159726 196188 159732 196200
rect 159784 196188 159790 196240
rect 161474 196188 161480 196240
rect 161532 196228 161538 196240
rect 162670 196228 162676 196240
rect 161532 196200 162676 196228
rect 161532 196188 161538 196200
rect 162670 196188 162676 196200
rect 162728 196188 162734 196240
rect 168742 196188 168748 196240
rect 168800 196228 168806 196240
rect 169570 196228 169576 196240
rect 168800 196200 169576 196228
rect 168800 196188 168806 196200
rect 169570 196188 169576 196200
rect 169628 196188 169634 196240
rect 138474 196160 138480 196172
rect 138032 196132 138480 196160
rect 137186 196052 137192 196104
rect 137244 196092 137250 196104
rect 137462 196092 137468 196104
rect 137244 196064 137468 196092
rect 137244 196052 137250 196064
rect 137462 196052 137468 196064
rect 137520 196052 137526 196104
rect 120166 195984 120172 196036
rect 120224 196024 120230 196036
rect 121454 196024 121460 196036
rect 120224 195996 121460 196024
rect 120224 195984 120230 195996
rect 121454 195984 121460 195996
rect 121512 195984 121518 196036
rect 134426 195916 134432 195968
rect 134484 195956 134490 195968
rect 135162 195956 135168 195968
rect 134484 195928 135168 195956
rect 134484 195916 134490 195928
rect 135162 195916 135168 195928
rect 135220 195916 135226 195968
rect 138032 195956 138060 196132
rect 138474 196120 138480 196132
rect 138532 196120 138538 196172
rect 153378 196120 153384 196172
rect 153436 196160 153442 196172
rect 153436 196132 153608 196160
rect 153436 196120 153442 196132
rect 153580 196104 153608 196132
rect 166166 196120 166172 196172
rect 166224 196160 166230 196172
rect 176194 196160 176200 196172
rect 166224 196132 176200 196160
rect 166224 196120 166230 196132
rect 176194 196120 176200 196132
rect 176252 196120 176258 196172
rect 138106 196052 138112 196104
rect 138164 196092 138170 196104
rect 139946 196092 139952 196104
rect 138164 196064 139952 196092
rect 138164 196052 138170 196064
rect 139946 196052 139952 196064
rect 140004 196052 140010 196104
rect 142338 196052 142344 196104
rect 142396 196092 142402 196104
rect 142798 196092 142804 196104
rect 142396 196064 142804 196092
rect 142396 196052 142402 196064
rect 142798 196052 142804 196064
rect 142856 196052 142862 196104
rect 153562 196052 153568 196104
rect 153620 196052 153626 196104
rect 161658 196052 161664 196104
rect 161716 196092 161722 196104
rect 162394 196092 162400 196104
rect 161716 196064 162400 196092
rect 161716 196052 161722 196064
rect 162394 196052 162400 196064
rect 162452 196052 162458 196104
rect 166994 196052 167000 196104
rect 167052 196092 167058 196104
rect 167362 196092 167368 196104
rect 167052 196064 167368 196092
rect 167052 196052 167058 196064
rect 167362 196052 167368 196064
rect 167420 196052 167426 196104
rect 173894 196052 173900 196104
rect 173952 196092 173958 196104
rect 174078 196092 174084 196104
rect 173952 196064 174084 196092
rect 173952 196052 173958 196064
rect 174078 196052 174084 196064
rect 174136 196052 174142 196104
rect 174170 196052 174176 196104
rect 174228 196092 174234 196104
rect 174814 196092 174820 196104
rect 174228 196064 174820 196092
rect 174228 196052 174234 196064
rect 174814 196052 174820 196064
rect 174872 196052 174878 196104
rect 148318 195984 148324 196036
rect 148376 196024 148382 196036
rect 148962 196024 148968 196036
rect 148376 195996 148968 196024
rect 148376 195984 148382 195996
rect 148962 195984 148968 195996
rect 149020 196024 149026 196036
rect 191190 196024 191196 196036
rect 149020 195996 191196 196024
rect 149020 195984 149026 195996
rect 191190 195984 191196 195996
rect 191248 195984 191254 196036
rect 215294 195984 215300 196036
rect 215352 196024 215358 196036
rect 215570 196024 215576 196036
rect 215352 195996 215576 196024
rect 215352 195984 215358 195996
rect 215570 195984 215576 195996
rect 215628 196024 215634 196036
rect 580350 196024 580356 196036
rect 215628 195996 580356 196024
rect 215628 195984 215634 195996
rect 580350 195984 580356 195996
rect 580408 195984 580414 196036
rect 138474 195956 138480 195968
rect 138032 195928 138480 195956
rect 138474 195916 138480 195928
rect 138532 195916 138538 195968
rect 139946 195916 139952 195968
rect 140004 195956 140010 195968
rect 140406 195956 140412 195968
rect 140004 195928 140412 195956
rect 140004 195916 140010 195928
rect 140406 195916 140412 195928
rect 140464 195916 140470 195968
rect 149606 195916 149612 195968
rect 149664 195956 149670 195968
rect 149882 195956 149888 195968
rect 149664 195928 149888 195956
rect 149664 195916 149670 195928
rect 149882 195916 149888 195928
rect 149940 195916 149946 195968
rect 156046 195916 156052 195968
rect 156104 195956 156110 195968
rect 157058 195956 157064 195968
rect 156104 195928 157064 195956
rect 156104 195916 156110 195928
rect 157058 195916 157064 195928
rect 157116 195916 157122 195968
rect 160462 195916 160468 195968
rect 160520 195956 160526 195968
rect 161290 195956 161296 195968
rect 160520 195928 161296 195956
rect 160520 195916 160526 195928
rect 161290 195916 161296 195928
rect 161348 195916 161354 195968
rect 163314 195916 163320 195968
rect 163372 195956 163378 195968
rect 193214 195956 193220 195968
rect 163372 195928 193220 195956
rect 163372 195916 163378 195928
rect 193214 195916 193220 195928
rect 193272 195956 193278 195968
rect 197446 195956 197452 195968
rect 193272 195928 197452 195956
rect 193272 195916 193278 195928
rect 197446 195916 197452 195928
rect 197504 195916 197510 195968
rect 108298 195848 108304 195900
rect 108356 195888 108362 195900
rect 171318 195888 171324 195900
rect 108356 195860 171324 195888
rect 108356 195848 108362 195860
rect 171318 195848 171324 195860
rect 171376 195888 171382 195900
rect 192938 195888 192944 195900
rect 171376 195860 192944 195888
rect 171376 195848 171382 195860
rect 192938 195848 192944 195860
rect 192996 195848 193002 195900
rect 108482 195780 108488 195832
rect 108540 195820 108546 195832
rect 174446 195820 174452 195832
rect 108540 195792 174452 195820
rect 108540 195780 108546 195792
rect 174446 195780 174452 195792
rect 174504 195820 174510 195832
rect 176286 195820 176292 195832
rect 174504 195792 176292 195820
rect 174504 195780 174510 195792
rect 176286 195780 176292 195792
rect 176344 195780 176350 195832
rect 108666 195712 108672 195764
rect 108724 195752 108730 195764
rect 170858 195752 170864 195764
rect 108724 195724 170864 195752
rect 108724 195712 108730 195724
rect 170858 195712 170864 195724
rect 170916 195752 170922 195764
rect 173894 195752 173900 195764
rect 170916 195724 173900 195752
rect 170916 195712 170922 195724
rect 173894 195712 173900 195724
rect 173952 195712 173958 195764
rect 198826 195712 198832 195764
rect 198884 195752 198890 195764
rect 212810 195752 212816 195764
rect 198884 195724 212816 195752
rect 198884 195712 198890 195724
rect 212810 195712 212816 195724
rect 212868 195752 212874 195764
rect 213822 195752 213828 195764
rect 212868 195724 213828 195752
rect 212868 195712 212874 195724
rect 213822 195712 213828 195724
rect 213880 195712 213886 195764
rect 117774 195644 117780 195696
rect 117832 195684 117838 195696
rect 147214 195684 147220 195696
rect 117832 195656 147220 195684
rect 117832 195644 117838 195656
rect 147214 195644 147220 195656
rect 147272 195644 147278 195696
rect 147766 195644 147772 195696
rect 147824 195684 147830 195696
rect 148502 195684 148508 195696
rect 147824 195656 148508 195684
rect 147824 195644 147830 195656
rect 148502 195644 148508 195656
rect 148560 195644 148566 195696
rect 154206 195644 154212 195696
rect 154264 195684 154270 195696
rect 154482 195684 154488 195696
rect 154264 195656 154488 195684
rect 154264 195644 154270 195656
rect 154482 195644 154488 195656
rect 154540 195644 154546 195696
rect 165430 195644 165436 195696
rect 165488 195684 165494 195696
rect 170766 195684 170772 195696
rect 165488 195656 170772 195684
rect 165488 195644 165494 195656
rect 170766 195644 170772 195656
rect 170824 195644 170830 195696
rect 174354 195644 174360 195696
rect 174412 195684 174418 195696
rect 174998 195684 175004 195696
rect 174412 195656 175004 195684
rect 174412 195644 174418 195656
rect 174998 195644 175004 195656
rect 175056 195684 175062 195696
rect 207290 195684 207296 195696
rect 175056 195656 207296 195684
rect 175056 195644 175062 195656
rect 207290 195644 207296 195656
rect 207348 195644 207354 195696
rect 122098 195576 122104 195628
rect 122156 195616 122162 195628
rect 148226 195616 148232 195628
rect 122156 195588 148232 195616
rect 122156 195576 122162 195588
rect 148226 195576 148232 195588
rect 148284 195576 148290 195628
rect 166350 195576 166356 195628
rect 166408 195616 166414 195628
rect 200298 195616 200304 195628
rect 166408 195588 200304 195616
rect 166408 195576 166414 195588
rect 200298 195576 200304 195588
rect 200356 195576 200362 195628
rect 117038 195508 117044 195560
rect 117096 195548 117102 195560
rect 149330 195548 149336 195560
rect 117096 195520 149336 195548
rect 117096 195508 117102 195520
rect 149330 195508 149336 195520
rect 149388 195508 149394 195560
rect 157242 195548 157248 195560
rect 151786 195520 157248 195548
rect 110230 195440 110236 195492
rect 110288 195480 110294 195492
rect 135530 195480 135536 195492
rect 110288 195452 135536 195480
rect 110288 195440 110294 195452
rect 135530 195440 135536 195452
rect 135588 195440 135594 195492
rect 137370 195440 137376 195492
rect 137428 195480 137434 195492
rect 137646 195480 137652 195492
rect 137428 195452 137652 195480
rect 137428 195440 137434 195452
rect 137646 195440 137652 195452
rect 137704 195440 137710 195492
rect 139394 195440 139400 195492
rect 139452 195480 139458 195492
rect 140406 195480 140412 195492
rect 139452 195452 140412 195480
rect 139452 195440 139458 195452
rect 140406 195440 140412 195452
rect 140464 195440 140470 195492
rect 100478 195372 100484 195424
rect 100536 195412 100542 195424
rect 133230 195412 133236 195424
rect 100536 195384 133236 195412
rect 100536 195372 100542 195384
rect 133230 195372 133236 195384
rect 133288 195372 133294 195424
rect 143994 195372 144000 195424
rect 144052 195412 144058 195424
rect 144178 195412 144184 195424
rect 144052 195384 144184 195412
rect 144052 195372 144058 195384
rect 144178 195372 144184 195384
rect 144236 195372 144242 195424
rect 109678 195304 109684 195356
rect 109736 195344 109742 195356
rect 151786 195344 151814 195520
rect 157242 195508 157248 195520
rect 157300 195508 157306 195560
rect 165706 195508 165712 195560
rect 165764 195548 165770 195560
rect 166534 195548 166540 195560
rect 165764 195520 166540 195548
rect 165764 195508 165770 195520
rect 166534 195508 166540 195520
rect 166592 195508 166598 195560
rect 168834 195508 168840 195560
rect 168892 195548 168898 195560
rect 170490 195548 170496 195560
rect 168892 195520 170496 195548
rect 168892 195508 168898 195520
rect 170490 195508 170496 195520
rect 170548 195508 170554 195560
rect 173066 195508 173072 195560
rect 173124 195548 173130 195560
rect 173526 195548 173532 195560
rect 173124 195520 173532 195548
rect 173124 195508 173130 195520
rect 173526 195508 173532 195520
rect 173584 195508 173590 195560
rect 179322 195508 179328 195560
rect 179380 195548 179386 195560
rect 215294 195548 215300 195560
rect 179380 195520 215300 195548
rect 179380 195508 179386 195520
rect 215294 195508 215300 195520
rect 215352 195508 215358 195560
rect 151998 195440 152004 195492
rect 152056 195480 152062 195492
rect 153010 195480 153016 195492
rect 152056 195452 153016 195480
rect 152056 195440 152062 195452
rect 153010 195440 153016 195452
rect 153068 195440 153074 195492
rect 164206 195452 166580 195480
rect 109736 195316 151814 195344
rect 109736 195304 109742 195316
rect 4798 195236 4804 195288
rect 4856 195276 4862 195288
rect 161750 195276 161756 195288
rect 4856 195248 161756 195276
rect 4856 195236 4862 195248
rect 161750 195236 161756 195248
rect 161808 195276 161814 195288
rect 164206 195276 164234 195452
rect 164878 195372 164884 195424
rect 164936 195412 164942 195424
rect 165154 195412 165160 195424
rect 164936 195384 165160 195412
rect 164936 195372 164942 195384
rect 165154 195372 165160 195384
rect 165212 195372 165218 195424
rect 165706 195372 165712 195424
rect 165764 195412 165770 195424
rect 166442 195412 166448 195424
rect 165764 195384 166448 195412
rect 165764 195372 165770 195384
rect 166442 195372 166448 195384
rect 166500 195372 166506 195424
rect 166552 195412 166580 195452
rect 178126 195440 178132 195492
rect 178184 195480 178190 195492
rect 215478 195480 215484 195492
rect 178184 195452 215484 195480
rect 178184 195440 178190 195452
rect 215478 195440 215484 195452
rect 215536 195440 215542 195492
rect 169662 195412 169668 195424
rect 166552 195384 169668 195412
rect 169662 195372 169668 195384
rect 169720 195372 169726 195424
rect 176286 195372 176292 195424
rect 176344 195412 176350 195424
rect 208578 195412 208584 195424
rect 176344 195384 208584 195412
rect 176344 195372 176350 195384
rect 208578 195372 208584 195384
rect 208636 195372 208642 195424
rect 214374 195372 214380 195424
rect 214432 195412 214438 195424
rect 323578 195412 323584 195424
rect 214432 195384 323584 195412
rect 214432 195372 214438 195384
rect 323578 195372 323584 195384
rect 323636 195372 323642 195424
rect 175458 195304 175464 195356
rect 175516 195344 175522 195356
rect 212534 195344 212540 195356
rect 175516 195316 212540 195344
rect 175516 195304 175522 195316
rect 212534 195304 212540 195316
rect 212592 195304 212598 195356
rect 213822 195304 213828 195356
rect 213880 195344 213886 195356
rect 574738 195344 574744 195356
rect 213880 195316 574744 195344
rect 213880 195304 213886 195316
rect 574738 195304 574744 195316
rect 574796 195304 574802 195356
rect 161808 195248 164234 195276
rect 161808 195236 161814 195248
rect 165154 195236 165160 195288
rect 165212 195276 165218 195288
rect 165338 195276 165344 195288
rect 165212 195248 165344 195276
rect 165212 195236 165218 195248
rect 165338 195236 165344 195248
rect 165396 195236 165402 195288
rect 165890 195236 165896 195288
rect 165948 195276 165954 195288
rect 166718 195276 166724 195288
rect 165948 195248 166724 195276
rect 165948 195236 165954 195248
rect 166718 195236 166724 195248
rect 166776 195236 166782 195288
rect 167362 195236 167368 195288
rect 167420 195276 167426 195288
rect 168282 195276 168288 195288
rect 167420 195248 168288 195276
rect 167420 195236 167426 195248
rect 168282 195236 168288 195248
rect 168340 195236 168346 195288
rect 169938 195236 169944 195288
rect 169996 195276 170002 195288
rect 209774 195276 209780 195288
rect 169996 195248 209780 195276
rect 169996 195236 170002 195248
rect 209774 195236 209780 195248
rect 209832 195276 209838 195288
rect 580810 195276 580816 195288
rect 209832 195248 580816 195276
rect 209832 195236 209838 195248
rect 580810 195236 580816 195248
rect 580868 195236 580874 195288
rect 108850 195168 108856 195220
rect 108908 195208 108914 195220
rect 108908 195180 122834 195208
rect 108908 195168 108914 195180
rect 122806 195004 122834 195180
rect 133322 195168 133328 195220
rect 133380 195208 133386 195220
rect 137922 195208 137928 195220
rect 133380 195180 137928 195208
rect 133380 195168 133386 195180
rect 137922 195168 137928 195180
rect 137980 195168 137986 195220
rect 178034 195208 178040 195220
rect 150084 195180 178040 195208
rect 130746 195100 130752 195152
rect 130804 195140 130810 195152
rect 139486 195140 139492 195152
rect 130804 195112 139492 195140
rect 130804 195100 130810 195112
rect 139486 195100 139492 195112
rect 139544 195100 139550 195152
rect 140958 195100 140964 195152
rect 141016 195140 141022 195152
rect 141326 195140 141332 195152
rect 141016 195112 141332 195140
rect 141016 195100 141022 195112
rect 141326 195100 141332 195112
rect 141384 195100 141390 195152
rect 145374 195100 145380 195152
rect 145432 195140 145438 195152
rect 150084 195140 150112 195180
rect 178034 195168 178040 195180
rect 178092 195168 178098 195220
rect 145432 195112 150112 195140
rect 145432 195100 145438 195112
rect 150986 195100 150992 195152
rect 151044 195140 151050 195152
rect 152734 195140 152740 195152
rect 151044 195112 152740 195140
rect 151044 195100 151050 195112
rect 152734 195100 152740 195112
rect 152792 195100 152798 195152
rect 158622 195100 158628 195152
rect 158680 195140 158686 195152
rect 182818 195140 182824 195152
rect 158680 195112 182824 195140
rect 158680 195100 158686 195112
rect 182818 195100 182824 195112
rect 182876 195100 182882 195152
rect 164602 195032 164608 195084
rect 164660 195072 164666 195084
rect 165522 195072 165528 195084
rect 164660 195044 165528 195072
rect 164660 195032 164666 195044
rect 165522 195032 165528 195044
rect 165580 195032 165586 195084
rect 169662 195032 169668 195084
rect 169720 195072 169726 195084
rect 180150 195072 180156 195084
rect 169720 195044 180156 195072
rect 169720 195032 169726 195044
rect 180150 195032 180156 195044
rect 180208 195032 180214 195084
rect 142522 195004 142528 195016
rect 122806 194976 142528 195004
rect 142522 194964 142528 194976
rect 142580 194964 142586 195016
rect 169938 194964 169944 195016
rect 169996 195004 170002 195016
rect 170674 195004 170680 195016
rect 169996 194976 170680 195004
rect 169996 194964 170002 194976
rect 170674 194964 170680 194976
rect 170732 194964 170738 195016
rect 173894 194964 173900 195016
rect 173952 195004 173958 195016
rect 174630 195004 174636 195016
rect 173952 194976 174636 195004
rect 173952 194964 173958 194976
rect 174630 194964 174636 194976
rect 174688 194964 174694 195016
rect 105722 194896 105728 194948
rect 105780 194936 105786 194948
rect 174354 194936 174360 194948
rect 105780 194908 122834 194936
rect 105780 194896 105786 194908
rect 122806 194868 122834 194908
rect 128326 194908 174360 194936
rect 128326 194868 128354 194908
rect 174354 194896 174360 194908
rect 174412 194896 174418 194948
rect 122806 194840 128354 194868
rect 141142 194828 141148 194880
rect 141200 194868 141206 194880
rect 141694 194868 141700 194880
rect 141200 194840 141700 194868
rect 141200 194828 141206 194840
rect 141694 194828 141700 194840
rect 141752 194828 141758 194880
rect 141878 194828 141884 194880
rect 141936 194868 141942 194880
rect 142522 194868 142528 194880
rect 141936 194840 142528 194868
rect 141936 194828 141942 194840
rect 142522 194828 142528 194840
rect 142580 194828 142586 194880
rect 165062 194828 165068 194880
rect 165120 194868 165126 194880
rect 165430 194868 165436 194880
rect 165120 194840 165436 194868
rect 165120 194828 165126 194840
rect 165430 194828 165436 194840
rect 165488 194828 165494 194880
rect 169018 194828 169024 194880
rect 169076 194868 169082 194880
rect 178770 194868 178776 194880
rect 169076 194840 178776 194868
rect 169076 194828 169082 194840
rect 178770 194828 178776 194840
rect 178828 194828 178834 194880
rect 128630 194760 128636 194812
rect 128688 194800 128694 194812
rect 132034 194800 132040 194812
rect 128688 194772 132040 194800
rect 128688 194760 128694 194772
rect 132034 194760 132040 194772
rect 132092 194760 132098 194812
rect 166534 194760 166540 194812
rect 166592 194800 166598 194812
rect 171870 194800 171876 194812
rect 166592 194772 171876 194800
rect 166592 194760 166598 194772
rect 171870 194760 171876 194772
rect 171928 194760 171934 194812
rect 133230 194692 133236 194744
rect 133288 194732 133294 194744
rect 141234 194732 141240 194744
rect 133288 194704 141240 194732
rect 133288 194692 133294 194704
rect 141234 194692 141240 194704
rect 141292 194692 141298 194744
rect 130654 194624 130660 194676
rect 130712 194664 130718 194676
rect 140038 194664 140044 194676
rect 130712 194636 140044 194664
rect 130712 194624 130718 194636
rect 140038 194624 140044 194636
rect 140096 194624 140102 194676
rect 202230 194624 202236 194676
rect 202288 194664 202294 194676
rect 214006 194664 214012 194676
rect 202288 194636 214012 194664
rect 202288 194624 202294 194636
rect 214006 194624 214012 194636
rect 214064 194664 214070 194676
rect 214374 194664 214380 194676
rect 214064 194636 214380 194664
rect 214064 194624 214070 194636
rect 214374 194624 214380 194636
rect 214432 194624 214438 194676
rect 96338 194556 96344 194608
rect 96396 194596 96402 194608
rect 103606 194596 103612 194608
rect 96396 194568 103612 194596
rect 96396 194556 96402 194568
rect 103606 194556 103612 194568
rect 103664 194596 103670 194608
rect 104618 194596 104624 194608
rect 103664 194568 104624 194596
rect 103664 194556 103670 194568
rect 104618 194556 104624 194568
rect 104676 194556 104682 194608
rect 178034 194556 178040 194608
rect 178092 194596 178098 194608
rect 580258 194596 580264 194608
rect 178092 194568 580264 194596
rect 178092 194556 178098 194568
rect 580258 194556 580264 194568
rect 580316 194556 580322 194608
rect 104342 194488 104348 194540
rect 104400 194528 104406 194540
rect 157426 194528 157432 194540
rect 104400 194500 157432 194528
rect 104400 194488 104406 194500
rect 157426 194488 157432 194500
rect 157484 194488 157490 194540
rect 163222 194488 163228 194540
rect 163280 194528 163286 194540
rect 163866 194528 163872 194540
rect 163280 194500 163872 194528
rect 163280 194488 163286 194500
rect 163866 194488 163872 194500
rect 163924 194488 163930 194540
rect 189994 194488 190000 194540
rect 190052 194528 190058 194540
rect 191834 194528 191840 194540
rect 190052 194500 191840 194528
rect 190052 194488 190058 194500
rect 191834 194488 191840 194500
rect 191892 194488 191898 194540
rect 107010 194420 107016 194472
rect 107068 194460 107074 194472
rect 114370 194460 114376 194472
rect 107068 194432 114376 194460
rect 107068 194420 107074 194432
rect 114370 194420 114376 194432
rect 114428 194420 114434 194472
rect 164786 194420 164792 194472
rect 164844 194460 164850 194472
rect 190914 194460 190920 194472
rect 164844 194432 190920 194460
rect 164844 194420 164850 194432
rect 190914 194420 190920 194432
rect 190972 194460 190978 194472
rect 202966 194460 202972 194472
rect 190972 194432 202972 194460
rect 190972 194420 190978 194432
rect 202966 194420 202972 194432
rect 203024 194420 203030 194472
rect 132218 194352 132224 194404
rect 132276 194392 132282 194404
rect 133414 194392 133420 194404
rect 132276 194364 133420 194392
rect 132276 194352 132282 194364
rect 133414 194352 133420 194364
rect 133472 194392 133478 194404
rect 207014 194392 207020 194404
rect 133472 194364 207020 194392
rect 133472 194352 133478 194364
rect 207014 194352 207020 194364
rect 207072 194352 207078 194404
rect 103146 194284 103152 194336
rect 103204 194324 103210 194336
rect 177114 194324 177120 194336
rect 103204 194296 177120 194324
rect 103204 194284 103210 194296
rect 177114 194284 177120 194296
rect 177172 194284 177178 194336
rect 195974 194284 195980 194336
rect 196032 194324 196038 194336
rect 204438 194324 204444 194336
rect 196032 194296 204444 194324
rect 196032 194284 196038 194296
rect 204438 194284 204444 194296
rect 204496 194284 204502 194336
rect 94590 194216 94596 194268
rect 94648 194256 94654 194268
rect 166994 194256 167000 194268
rect 94648 194228 167000 194256
rect 94648 194216 94654 194228
rect 166994 194216 167000 194228
rect 167052 194216 167058 194268
rect 170398 194216 170404 194268
rect 170456 194256 170462 194268
rect 189626 194256 189632 194268
rect 170456 194228 189632 194256
rect 170456 194216 170462 194228
rect 189626 194216 189632 194228
rect 189684 194256 189690 194268
rect 189994 194256 190000 194268
rect 189684 194228 190000 194256
rect 189684 194216 189690 194228
rect 189994 194216 190000 194228
rect 190052 194216 190058 194268
rect 103054 194148 103060 194200
rect 103112 194188 103118 194200
rect 176010 194188 176016 194200
rect 103112 194160 176016 194188
rect 103112 194148 103118 194160
rect 176010 194148 176016 194160
rect 176068 194188 176074 194200
rect 176068 194160 180794 194188
rect 176068 194148 176074 194160
rect 104618 194080 104624 194132
rect 104676 194120 104682 194132
rect 114738 194120 114744 194132
rect 104676 194092 114744 194120
rect 104676 194080 104682 194092
rect 114738 194080 114744 194092
rect 114796 194080 114802 194132
rect 118050 194080 118056 194132
rect 118108 194120 118114 194132
rect 121362 194120 121368 194132
rect 118108 194092 121368 194120
rect 118108 194080 118114 194092
rect 121362 194080 121368 194092
rect 121420 194120 121426 194132
rect 153194 194120 153200 194132
rect 121420 194092 153200 194120
rect 121420 194080 121426 194092
rect 153194 194080 153200 194092
rect 153252 194080 153258 194132
rect 180766 194120 180794 194160
rect 190086 194148 190092 194200
rect 190144 194188 190150 194200
rect 205634 194188 205640 194200
rect 190144 194160 205640 194188
rect 190144 194148 190150 194160
rect 205634 194148 205640 194160
rect 205692 194148 205698 194200
rect 200482 194120 200488 194132
rect 180766 194092 200488 194120
rect 200482 194080 200488 194092
rect 200540 194080 200546 194132
rect 114370 194012 114376 194064
rect 114428 194052 114434 194064
rect 146202 194052 146208 194064
rect 114428 194024 146208 194052
rect 114428 194012 114434 194024
rect 146202 194012 146208 194024
rect 146260 194012 146266 194064
rect 157610 194012 157616 194064
rect 157668 194052 157674 194064
rect 174538 194052 174544 194064
rect 157668 194024 174544 194052
rect 157668 194012 157674 194024
rect 174538 194012 174544 194024
rect 174596 194012 174602 194064
rect 177114 194012 177120 194064
rect 177172 194052 177178 194064
rect 177850 194052 177856 194064
rect 177172 194024 177856 194052
rect 177172 194012 177178 194024
rect 177850 194012 177856 194024
rect 177908 194052 177914 194064
rect 203058 194052 203064 194064
rect 177908 194024 203064 194052
rect 177908 194012 177914 194024
rect 203058 194012 203064 194024
rect 203116 194012 203122 194064
rect 102594 193944 102600 193996
rect 102652 193984 102658 193996
rect 126974 193984 126980 193996
rect 102652 193956 126980 193984
rect 102652 193944 102658 193956
rect 126974 193944 126980 193956
rect 127032 193944 127038 193996
rect 149330 193944 149336 193996
rect 149388 193984 149394 193996
rect 149974 193984 149980 193996
rect 149388 193956 149980 193984
rect 149388 193944 149394 193956
rect 149974 193944 149980 193956
rect 150032 193944 150038 193996
rect 157978 193944 157984 193996
rect 158036 193984 158042 193996
rect 196618 193984 196624 193996
rect 158036 193956 196624 193984
rect 158036 193944 158042 193956
rect 196618 193944 196624 193956
rect 196676 193944 196682 193996
rect 198826 193944 198832 193996
rect 198884 193984 198890 193996
rect 502978 193984 502984 193996
rect 198884 193956 502984 193984
rect 198884 193944 198890 193956
rect 502978 193944 502984 193956
rect 503036 193944 503042 193996
rect 94590 193876 94596 193928
rect 94648 193916 94654 193928
rect 103514 193916 103520 193928
rect 94648 193888 103520 193916
rect 94648 193876 94654 193888
rect 103514 193876 103520 193888
rect 103572 193916 103578 193928
rect 104342 193916 104348 193928
rect 103572 193888 104348 193916
rect 103572 193876 103578 193888
rect 104342 193876 104348 193888
rect 104400 193876 104406 193928
rect 104618 193876 104624 193928
rect 104676 193916 104682 193928
rect 137094 193916 137100 193928
rect 104676 193888 137100 193916
rect 104676 193876 104682 193888
rect 137094 193876 137100 193888
rect 137152 193876 137158 193928
rect 146202 193876 146208 193928
rect 146260 193916 146266 193928
rect 151814 193916 151820 193928
rect 146260 193888 151820 193916
rect 146260 193876 146266 193888
rect 151814 193876 151820 193888
rect 151872 193876 151878 193928
rect 162578 193876 162584 193928
rect 162636 193916 162642 193928
rect 195974 193916 195980 193928
rect 162636 193888 195980 193916
rect 162636 193876 162642 193888
rect 195974 193876 195980 193888
rect 196032 193916 196038 193928
rect 580626 193916 580632 193928
rect 196032 193888 580632 193916
rect 196032 193876 196038 193888
rect 580626 193876 580632 193888
rect 580684 193876 580690 193928
rect 3418 193808 3424 193860
rect 3476 193848 3482 193860
rect 114094 193848 114100 193860
rect 3476 193820 114100 193848
rect 3476 193808 3482 193820
rect 114094 193808 114100 193820
rect 114152 193848 114158 193860
rect 146662 193848 146668 193860
rect 114152 193820 146668 193848
rect 114152 193808 114158 193820
rect 146662 193808 146668 193820
rect 146720 193808 146726 193860
rect 120350 193740 120356 193792
rect 120408 193780 120414 193792
rect 142062 193780 142068 193792
rect 120408 193752 142068 193780
rect 120408 193740 120414 193752
rect 142062 193740 142068 193752
rect 142120 193740 142126 193792
rect 171502 193740 171508 193792
rect 171560 193780 171566 193792
rect 188614 193780 188620 193792
rect 171560 193752 188620 193780
rect 171560 193740 171566 193752
rect 188614 193740 188620 193752
rect 188672 193740 188678 193792
rect 122006 193672 122012 193724
rect 122064 193712 122070 193724
rect 135806 193712 135812 193724
rect 122064 193684 135812 193712
rect 122064 193672 122070 193684
rect 135806 193672 135812 193684
rect 135864 193672 135870 193724
rect 165614 193672 165620 193724
rect 165672 193712 165678 193724
rect 185578 193712 185584 193724
rect 165672 193684 185584 193712
rect 165672 193672 165678 193684
rect 185578 193672 185584 193684
rect 185636 193672 185642 193724
rect 152458 193604 152464 193656
rect 152516 193644 152522 193656
rect 328454 193644 328460 193656
rect 152516 193616 328460 193644
rect 152516 193604 152522 193616
rect 328454 193604 328460 193616
rect 328512 193604 328518 193656
rect 148502 193536 148508 193588
rect 148560 193576 148566 193588
rect 579798 193576 579804 193588
rect 148560 193548 579804 193576
rect 148560 193536 148566 193548
rect 579798 193536 579804 193548
rect 579856 193536 579862 193588
rect 90450 193468 90456 193520
rect 90508 193508 90514 193520
rect 164878 193508 164884 193520
rect 90508 193480 164884 193508
rect 90508 193468 90514 193480
rect 164878 193468 164884 193480
rect 164936 193468 164942 193520
rect 164970 193468 164976 193520
rect 165028 193508 165034 193520
rect 165614 193508 165620 193520
rect 165028 193480 165620 193508
rect 165028 193468 165034 193480
rect 165614 193468 165620 193480
rect 165672 193468 165678 193520
rect 114922 193400 114928 193452
rect 114980 193440 114986 193452
rect 147674 193440 147680 193452
rect 114980 193412 147680 193440
rect 114980 193400 114986 193412
rect 147674 193400 147680 193412
rect 147732 193400 147738 193452
rect 157794 193400 157800 193452
rect 157852 193440 157858 193452
rect 158346 193440 158352 193452
rect 157852 193412 158352 193440
rect 157852 193400 157858 193412
rect 158346 193400 158352 193412
rect 158404 193400 158410 193452
rect 178034 193332 178040 193384
rect 178092 193372 178098 193384
rect 178862 193372 178868 193384
rect 178092 193344 178868 193372
rect 178092 193332 178098 193344
rect 178862 193332 178868 193344
rect 178920 193332 178926 193384
rect 96614 193264 96620 193316
rect 96672 193304 96678 193316
rect 118694 193304 118700 193316
rect 96672 193276 118700 193304
rect 96672 193264 96678 193276
rect 118694 193264 118700 193276
rect 118752 193264 118758 193316
rect 104158 193196 104164 193248
rect 104216 193236 104222 193248
rect 112806 193236 112812 193248
rect 104216 193208 112812 193236
rect 104216 193196 104222 193208
rect 112806 193196 112812 193208
rect 112864 193236 112870 193248
rect 112864 193208 113174 193236
rect 112864 193196 112870 193208
rect 113146 193100 113174 193208
rect 124950 193196 124956 193248
rect 125008 193236 125014 193248
rect 132310 193236 132316 193248
rect 125008 193208 132316 193236
rect 125008 193196 125014 193208
rect 132310 193196 132316 193208
rect 132368 193196 132374 193248
rect 134518 193196 134524 193248
rect 134576 193236 134582 193248
rect 134576 193208 135300 193236
rect 134576 193196 134582 193208
rect 135272 193168 135300 193208
rect 170490 193196 170496 193248
rect 170548 193236 170554 193248
rect 188706 193236 188712 193248
rect 170548 193208 188712 193236
rect 170548 193196 170554 193208
rect 188706 193196 188712 193208
rect 188764 193196 188770 193248
rect 142154 193168 142160 193180
rect 135272 193140 142160 193168
rect 142154 193128 142160 193140
rect 142212 193168 142218 193180
rect 580442 193168 580448 193180
rect 142212 193140 580448 193168
rect 142212 193128 142218 193140
rect 580442 193128 580448 193140
rect 580500 193128 580506 193180
rect 138014 193100 138020 193112
rect 113146 193072 138020 193100
rect 138014 193060 138020 193072
rect 138072 193060 138078 193112
rect 140038 193060 140044 193112
rect 140096 193100 140102 193112
rect 142982 193100 142988 193112
rect 140096 193072 142988 193100
rect 140096 193060 140102 193072
rect 142982 193060 142988 193072
rect 143040 193100 143046 193112
rect 576394 193100 576400 193112
rect 143040 193072 576400 193100
rect 143040 193060 143046 193072
rect 576394 193060 576400 193072
rect 576452 193060 576458 193112
rect 132310 192992 132316 193044
rect 132368 193032 132374 193044
rect 145742 193032 145748 193044
rect 132368 193004 145748 193032
rect 132368 192992 132374 193004
rect 145742 192992 145748 193004
rect 145800 193032 145806 193044
rect 577590 193032 577596 193044
rect 145800 193004 577596 193032
rect 145800 192992 145806 193004
rect 577590 192992 577596 193004
rect 577648 192992 577654 193044
rect 132954 192924 132960 192976
rect 133012 192964 133018 192976
rect 201494 192964 201500 192976
rect 133012 192936 201500 192964
rect 133012 192924 133018 192936
rect 201494 192924 201500 192936
rect 201552 192924 201558 192976
rect 109862 192856 109868 192908
rect 109920 192896 109926 192908
rect 163682 192896 163688 192908
rect 109920 192868 163688 192896
rect 109920 192856 109926 192868
rect 163682 192856 163688 192868
rect 163740 192856 163746 192908
rect 172238 192856 172244 192908
rect 172296 192896 172302 192908
rect 172296 192868 190454 192896
rect 172296 192856 172302 192868
rect 108114 192788 108120 192840
rect 108172 192828 108178 192840
rect 138198 192828 138204 192840
rect 108172 192800 138204 192828
rect 108172 192788 108178 192800
rect 138198 192788 138204 192800
rect 138256 192788 138262 192840
rect 147674 192788 147680 192840
rect 147732 192828 147738 192840
rect 148686 192828 148692 192840
rect 147732 192800 148692 192828
rect 147732 192788 147738 192800
rect 148686 192788 148692 192800
rect 148744 192828 148750 192840
rect 189442 192828 189448 192840
rect 148744 192800 189448 192828
rect 148744 192788 148750 192800
rect 189442 192788 189448 192800
rect 189500 192788 189506 192840
rect 190426 192828 190454 192868
rect 194686 192828 194692 192840
rect 190426 192800 194692 192828
rect 194686 192788 194692 192800
rect 194744 192828 194750 192840
rect 204714 192828 204720 192840
rect 194744 192800 204720 192828
rect 194744 192788 194750 192800
rect 204714 192788 204720 192800
rect 204772 192788 204778 192840
rect 113082 192720 113088 192772
rect 113140 192760 113146 192772
rect 146294 192760 146300 192772
rect 113140 192732 146300 192760
rect 113140 192720 113146 192732
rect 146294 192720 146300 192732
rect 146352 192720 146358 192772
rect 152182 192720 152188 192772
rect 152240 192760 152246 192772
rect 152734 192760 152740 192772
rect 152240 192732 152740 192760
rect 152240 192720 152246 192732
rect 152734 192720 152740 192732
rect 152792 192720 152798 192772
rect 174262 192720 174268 192772
rect 174320 192760 174326 192772
rect 208394 192760 208400 192772
rect 174320 192732 208400 192760
rect 174320 192720 174326 192732
rect 208394 192720 208400 192732
rect 208452 192720 208458 192772
rect 103330 192652 103336 192704
rect 103388 192692 103394 192704
rect 135438 192692 135444 192704
rect 103388 192664 135444 192692
rect 103388 192652 103394 192664
rect 135438 192652 135444 192664
rect 135496 192652 135502 192704
rect 142430 192652 142436 192704
rect 142488 192692 142494 192704
rect 332594 192692 332600 192704
rect 142488 192664 332600 192692
rect 142488 192652 142494 192664
rect 332594 192652 332600 192664
rect 332652 192652 332658 192704
rect 93302 192584 93308 192636
rect 93360 192624 93366 192636
rect 101858 192624 101864 192636
rect 93360 192596 101864 192624
rect 93360 192584 93366 192596
rect 101858 192584 101864 192596
rect 101916 192624 101922 192636
rect 136358 192624 136364 192636
rect 101916 192596 136364 192624
rect 101916 192584 101922 192596
rect 136358 192584 136364 192596
rect 136416 192584 136422 192636
rect 171686 192584 171692 192636
rect 171744 192624 171750 192636
rect 217134 192624 217140 192636
rect 171744 192596 217140 192624
rect 171744 192584 171750 192596
rect 217134 192584 217140 192596
rect 217192 192624 217198 192636
rect 561122 192624 561128 192636
rect 217192 192596 561128 192624
rect 217192 192584 217198 192596
rect 561122 192584 561128 192596
rect 561180 192584 561186 192636
rect 86218 192516 86224 192568
rect 86276 192556 86282 192568
rect 99006 192556 99012 192568
rect 86276 192528 99012 192556
rect 86276 192516 86282 192528
rect 99006 192516 99012 192528
rect 99064 192556 99070 192568
rect 128630 192556 128636 192568
rect 99064 192528 128636 192556
rect 99064 192516 99070 192528
rect 128630 192516 128636 192528
rect 128688 192516 128694 192568
rect 132310 192516 132316 192568
rect 132368 192556 132374 192568
rect 132954 192556 132960 192568
rect 132368 192528 132960 192556
rect 132368 192516 132374 192528
rect 132954 192516 132960 192528
rect 133012 192516 133018 192568
rect 160830 192516 160836 192568
rect 160888 192556 160894 192568
rect 173250 192556 173256 192568
rect 160888 192528 173256 192556
rect 160888 192516 160894 192528
rect 173250 192516 173256 192528
rect 173308 192516 173314 192568
rect 175090 192516 175096 192568
rect 175148 192556 175154 192568
rect 214282 192556 214288 192568
rect 175148 192528 214288 192556
rect 175148 192516 175154 192528
rect 214282 192516 214288 192528
rect 214340 192556 214346 192568
rect 580902 192556 580908 192568
rect 214340 192528 580908 192556
rect 214340 192516 214346 192528
rect 580902 192516 580908 192528
rect 580960 192516 580966 192568
rect 3418 192448 3424 192500
rect 3476 192488 3482 192500
rect 124214 192488 124220 192500
rect 3476 192460 124220 192488
rect 3476 192448 3482 192460
rect 124214 192448 124220 192460
rect 124272 192488 124278 192500
rect 125502 192488 125508 192500
rect 124272 192460 125508 192488
rect 124272 192448 124278 192460
rect 125502 192448 125508 192460
rect 125560 192448 125566 192500
rect 127618 192448 127624 192500
rect 127676 192488 127682 192500
rect 147214 192488 147220 192500
rect 127676 192460 147220 192488
rect 127676 192448 127682 192460
rect 147214 192448 147220 192460
rect 147272 192448 147278 192500
rect 156782 192448 156788 192500
rect 156840 192488 156846 192500
rect 197354 192488 197360 192500
rect 156840 192460 197360 192488
rect 156840 192448 156846 192460
rect 197354 192448 197360 192460
rect 197412 192448 197418 192500
rect 208394 192448 208400 192500
rect 208452 192488 208458 192500
rect 208946 192488 208952 192500
rect 208452 192460 208952 192488
rect 208452 192448 208458 192460
rect 208946 192448 208952 192460
rect 209004 192488 209010 192500
rect 577866 192488 577872 192500
rect 209004 192460 577872 192488
rect 209004 192448 209010 192460
rect 577866 192448 577872 192460
rect 577924 192448 577930 192500
rect 116394 192380 116400 192432
rect 116452 192420 116458 192432
rect 139762 192420 139768 192432
rect 116452 192392 139768 192420
rect 116452 192380 116458 192392
rect 139762 192380 139768 192392
rect 139820 192380 139826 192432
rect 175182 192380 175188 192432
rect 175240 192420 175246 192432
rect 189718 192420 189724 192432
rect 175240 192392 189724 192420
rect 175240 192380 175246 192392
rect 189718 192380 189724 192392
rect 189776 192380 189782 192432
rect 118694 192312 118700 192364
rect 118752 192352 118758 192364
rect 144086 192352 144092 192364
rect 118752 192324 144092 192352
rect 118752 192312 118758 192324
rect 144086 192312 144092 192324
rect 144144 192312 144150 192364
rect 114738 192244 114744 192296
rect 114796 192284 114802 192296
rect 144822 192284 144828 192296
rect 114796 192256 144828 192284
rect 114796 192244 114802 192256
rect 144822 192244 144828 192256
rect 144880 192244 144886 192296
rect 109402 192176 109408 192228
rect 109460 192216 109466 192228
rect 140038 192216 140044 192228
rect 109460 192188 140044 192216
rect 109460 192176 109466 192188
rect 140038 192176 140044 192188
rect 140096 192176 140102 192228
rect 101766 191836 101772 191888
rect 101824 191876 101830 191888
rect 105630 191876 105636 191888
rect 101824 191848 105636 191876
rect 101824 191836 101830 191848
rect 105630 191836 105636 191848
rect 105688 191836 105694 191888
rect 100202 191768 100208 191820
rect 100260 191808 100266 191820
rect 111978 191808 111984 191820
rect 100260 191780 111984 191808
rect 100260 191768 100266 191780
rect 111978 191768 111984 191780
rect 112036 191768 112042 191820
rect 136910 191768 136916 191820
rect 136968 191808 136974 191820
rect 137646 191808 137652 191820
rect 136968 191780 137652 191808
rect 136968 191768 136974 191780
rect 137646 191768 137652 191780
rect 137704 191768 137710 191820
rect 141510 191768 141516 191820
rect 141568 191808 141574 191820
rect 144270 191808 144276 191820
rect 141568 191780 144276 191808
rect 141568 191768 141574 191780
rect 144270 191768 144276 191780
rect 144328 191808 144334 191820
rect 579154 191808 579160 191820
rect 144328 191780 579160 191808
rect 144328 191768 144334 191780
rect 579154 191768 579160 191780
rect 579212 191768 579218 191820
rect 103238 191700 103244 191752
rect 103296 191740 103302 191752
rect 134426 191740 134432 191752
rect 103296 191712 134432 191740
rect 103296 191700 103302 191712
rect 134426 191700 134432 191712
rect 134484 191700 134490 191752
rect 137186 191700 137192 191752
rect 137244 191740 137250 191752
rect 137922 191740 137928 191752
rect 137244 191712 137928 191740
rect 137244 191700 137250 191712
rect 137922 191700 137928 191712
rect 137980 191700 137986 191752
rect 139394 191700 139400 191752
rect 139452 191740 139458 191752
rect 140682 191740 140688 191752
rect 139452 191712 140688 191740
rect 139452 191700 139458 191712
rect 140682 191700 140688 191712
rect 140740 191740 140746 191752
rect 256694 191740 256700 191752
rect 140740 191712 256700 191740
rect 140740 191700 140746 191712
rect 256694 191700 256700 191712
rect 256752 191700 256758 191752
rect 93118 191632 93124 191684
rect 93176 191672 93182 191684
rect 165430 191672 165436 191684
rect 93176 191644 165436 191672
rect 93176 191632 93182 191644
rect 165430 191632 165436 191644
rect 165488 191632 165494 191684
rect 102686 191564 102692 191616
rect 102744 191604 102750 191616
rect 172606 191604 172612 191616
rect 102744 191576 172612 191604
rect 102744 191564 102750 191576
rect 172606 191564 172612 191576
rect 172664 191604 172670 191616
rect 188798 191604 188804 191616
rect 172664 191576 188804 191604
rect 172664 191564 172670 191576
rect 188798 191564 188804 191576
rect 188856 191564 188862 191616
rect 97442 191496 97448 191548
rect 97500 191536 97506 191548
rect 111150 191536 111156 191548
rect 97500 191508 111156 191536
rect 97500 191496 97506 191508
rect 111150 191496 111156 191508
rect 111208 191496 111214 191548
rect 117222 191496 117228 191548
rect 117280 191536 117286 191548
rect 161934 191536 161940 191548
rect 117280 191508 161940 191536
rect 117280 191496 117286 191508
rect 161934 191496 161940 191508
rect 161992 191536 161998 191548
rect 162670 191536 162676 191548
rect 161992 191508 162676 191536
rect 161992 191496 161998 191508
rect 162670 191496 162676 191508
rect 162728 191496 162734 191548
rect 176102 191496 176108 191548
rect 176160 191536 176166 191548
rect 200850 191536 200856 191548
rect 176160 191508 200856 191536
rect 176160 191496 176166 191508
rect 200850 191496 200856 191508
rect 200908 191496 200914 191548
rect 97258 191428 97264 191480
rect 97316 191468 97322 191480
rect 108666 191468 108672 191480
rect 97316 191440 108672 191468
rect 97316 191428 97322 191440
rect 108666 191428 108672 191440
rect 108724 191468 108730 191480
rect 142246 191468 142252 191480
rect 108724 191440 142252 191468
rect 108724 191428 108730 191440
rect 142246 191428 142252 191440
rect 142304 191428 142310 191480
rect 159634 191428 159640 191480
rect 159692 191468 159698 191480
rect 185670 191468 185676 191480
rect 159692 191440 185676 191468
rect 159692 191428 159698 191440
rect 185670 191428 185676 191440
rect 185728 191428 185734 191480
rect 100202 191360 100208 191412
rect 100260 191400 100266 191412
rect 133874 191400 133880 191412
rect 100260 191372 133880 191400
rect 100260 191360 100266 191372
rect 133874 191360 133880 191372
rect 133932 191360 133938 191412
rect 135530 191360 135536 191412
rect 135588 191400 135594 191412
rect 136542 191400 136548 191412
rect 135588 191372 136548 191400
rect 135588 191360 135594 191372
rect 136542 191360 136548 191372
rect 136600 191360 136606 191412
rect 137094 191360 137100 191412
rect 137152 191400 137158 191412
rect 137738 191400 137744 191412
rect 137152 191372 137744 191400
rect 137152 191360 137158 191372
rect 137738 191360 137744 191372
rect 137796 191360 137802 191412
rect 155310 191360 155316 191412
rect 155368 191400 155374 191412
rect 186406 191400 186412 191412
rect 155368 191372 186412 191400
rect 155368 191360 155374 191372
rect 186406 191360 186412 191372
rect 186464 191360 186470 191412
rect 100110 191292 100116 191344
rect 100168 191332 100174 191344
rect 117222 191332 117228 191344
rect 100168 191304 117228 191332
rect 100168 191292 100174 191304
rect 117222 191292 117228 191304
rect 117280 191332 117286 191344
rect 154482 191332 154488 191344
rect 117280 191304 154488 191332
rect 117280 191292 117286 191304
rect 154482 191292 154488 191304
rect 154540 191292 154546 191344
rect 162670 191292 162676 191344
rect 162728 191332 162734 191344
rect 196158 191332 196164 191344
rect 162728 191304 196164 191332
rect 162728 191292 162734 191304
rect 196158 191292 196164 191304
rect 196216 191292 196222 191344
rect 94682 191224 94688 191276
rect 94740 191264 94746 191276
rect 111794 191264 111800 191276
rect 94740 191236 111800 191264
rect 94740 191224 94746 191236
rect 111794 191224 111800 191236
rect 111852 191224 111858 191276
rect 115290 191224 115296 191276
rect 115348 191264 115354 191276
rect 150342 191264 150348 191276
rect 115348 191236 150348 191264
rect 115348 191224 115354 191236
rect 150342 191224 150348 191236
rect 150400 191224 150406 191276
rect 193950 191264 193956 191276
rect 153396 191236 193956 191264
rect 80054 191156 80060 191208
rect 80112 191196 80118 191208
rect 118602 191196 118608 191208
rect 80112 191168 118608 191196
rect 80112 191156 80118 191168
rect 118602 191156 118608 191168
rect 118660 191196 118666 191208
rect 153286 191196 153292 191208
rect 118660 191168 153292 191196
rect 118660 191156 118666 191168
rect 153286 191156 153292 191168
rect 153344 191156 153350 191208
rect 99098 191088 99104 191140
rect 99156 191128 99162 191140
rect 139394 191128 139400 191140
rect 99156 191100 139400 191128
rect 99156 191088 99162 191100
rect 139394 191088 139400 191100
rect 139452 191088 139458 191140
rect 109770 191020 109776 191072
rect 109828 191060 109834 191072
rect 119430 191060 119436 191072
rect 109828 191032 119436 191060
rect 109828 191020 109834 191032
rect 119430 191020 119436 191032
rect 119488 191060 119494 191072
rect 149054 191060 149060 191072
rect 119488 191032 149060 191060
rect 119488 191020 119494 191032
rect 149054 191020 149060 191032
rect 149112 191020 149118 191072
rect 107102 190952 107108 191004
rect 107160 190992 107166 191004
rect 115290 190992 115296 191004
rect 107160 190964 115296 190992
rect 107160 190952 107166 190964
rect 115290 190952 115296 190964
rect 115348 190952 115354 191004
rect 132678 190952 132684 191004
rect 132736 190992 132742 191004
rect 132862 190992 132868 191004
rect 132736 190964 132868 190992
rect 132736 190952 132742 190964
rect 132862 190952 132868 190964
rect 132920 190952 132926 191004
rect 134058 190952 134064 191004
rect 134116 190992 134122 191004
rect 134794 190992 134800 191004
rect 134116 190964 134800 190992
rect 134116 190952 134122 190964
rect 134794 190952 134800 190964
rect 134852 190952 134858 191004
rect 135714 190952 135720 191004
rect 135772 190992 135778 191004
rect 136450 190992 136456 191004
rect 135772 190964 136456 190992
rect 135772 190952 135778 190964
rect 136450 190952 136456 190964
rect 136508 190952 136514 191004
rect 115842 190884 115848 190936
rect 115900 190924 115906 190936
rect 152090 190924 152096 190936
rect 115900 190896 137784 190924
rect 115900 190884 115906 190896
rect 132678 190816 132684 190868
rect 132736 190856 132742 190868
rect 133414 190856 133420 190868
rect 132736 190828 133420 190856
rect 132736 190816 132742 190828
rect 133414 190816 133420 190828
rect 133472 190816 133478 190868
rect 137002 190816 137008 190868
rect 137060 190856 137066 190868
rect 137554 190856 137560 190868
rect 137060 190828 137560 190856
rect 137060 190816 137066 190828
rect 137554 190816 137560 190828
rect 137612 190816 137618 190868
rect 137756 190856 137784 190896
rect 137940 190896 152096 190924
rect 137940 190856 137968 190896
rect 152090 190884 152096 190896
rect 152148 190924 152154 190936
rect 153396 190924 153424 191236
rect 193950 191224 193956 191236
rect 194008 191224 194014 191276
rect 166994 191156 167000 191208
rect 167052 191196 167058 191208
rect 209130 191196 209136 191208
rect 167052 191168 209136 191196
rect 167052 191156 167058 191168
rect 209130 191156 209136 191168
rect 209188 191156 209194 191208
rect 159910 191088 159916 191140
rect 159968 191128 159974 191140
rect 183462 191128 183468 191140
rect 159968 191100 183468 191128
rect 159968 191088 159974 191100
rect 183462 191088 183468 191100
rect 183520 191128 183526 191140
rect 578878 191128 578884 191140
rect 183520 191100 578884 191128
rect 183520 191088 183526 191100
rect 578878 191088 578884 191100
rect 578936 191088 578942 191140
rect 155402 191020 155408 191072
rect 155460 191060 155466 191072
rect 155862 191060 155868 191072
rect 155460 191032 155868 191060
rect 155460 191020 155466 191032
rect 155862 191020 155868 191032
rect 155920 191020 155926 191072
rect 167270 190952 167276 191004
rect 167328 190992 167334 191004
rect 167546 190992 167552 191004
rect 167328 190964 167552 190992
rect 167328 190952 167334 190964
rect 167546 190952 167552 190964
rect 167604 190952 167610 191004
rect 152148 190896 153424 190924
rect 152148 190884 152154 190896
rect 137756 190828 137968 190856
rect 136910 190748 136916 190800
rect 136968 190788 136974 190800
rect 137370 190788 137376 190800
rect 136968 190760 137376 190788
rect 136968 190748 136974 190760
rect 137370 190748 137376 190760
rect 137428 190748 137434 190800
rect 130470 190680 130476 190732
rect 130528 190720 130534 190732
rect 141510 190720 141516 190732
rect 130528 190692 141516 190720
rect 130528 190680 130534 190692
rect 141510 190680 141516 190692
rect 141568 190680 141574 190732
rect 137186 190612 137192 190664
rect 137244 190652 137250 190664
rect 137830 190652 137836 190664
rect 137244 190624 137836 190652
rect 137244 190612 137250 190624
rect 137830 190612 137836 190624
rect 137888 190612 137894 190664
rect 8938 190476 8944 190528
rect 8996 190516 9002 190528
rect 100202 190516 100208 190528
rect 8996 190488 100208 190516
rect 8996 190476 9002 190488
rect 100202 190476 100208 190488
rect 100260 190476 100266 190528
rect 108574 190476 108580 190528
rect 108632 190516 108638 190528
rect 113174 190516 113180 190528
rect 108632 190488 113180 190516
rect 108632 190476 108638 190488
rect 113174 190476 113180 190488
rect 113232 190476 113238 190528
rect 168834 190476 168840 190528
rect 168892 190516 168898 190528
rect 199194 190516 199200 190528
rect 168892 190488 199200 190516
rect 168892 190476 168898 190488
rect 199194 190476 199200 190488
rect 199252 190476 199258 190528
rect 136634 190408 136640 190460
rect 136692 190448 136698 190460
rect 137278 190448 137284 190460
rect 136692 190420 137284 190448
rect 136692 190408 136698 190420
rect 137278 190408 137284 190420
rect 137336 190448 137342 190460
rect 582742 190448 582748 190460
rect 137336 190420 582748 190448
rect 137336 190408 137342 190420
rect 582742 190408 582748 190420
rect 582800 190408 582806 190460
rect 133230 190340 133236 190392
rect 133288 190380 133294 190392
rect 153102 190380 153108 190392
rect 133288 190352 153108 190380
rect 133288 190340 133294 190352
rect 153102 190340 153108 190352
rect 153160 190380 153166 190392
rect 577682 190380 577688 190392
rect 153160 190352 577688 190380
rect 153160 190340 153166 190352
rect 577682 190340 577688 190352
rect 577740 190340 577746 190392
rect 91738 190272 91744 190324
rect 91796 190312 91802 190324
rect 170490 190312 170496 190324
rect 91796 190284 170496 190312
rect 91796 190272 91802 190284
rect 170490 190272 170496 190284
rect 170548 190272 170554 190324
rect 171778 190272 171784 190324
rect 171836 190312 171842 190324
rect 191006 190312 191012 190324
rect 171836 190284 191012 190312
rect 171836 190272 171842 190284
rect 191006 190272 191012 190284
rect 191064 190272 191070 190324
rect 111794 190204 111800 190256
rect 111852 190244 111858 190256
rect 112714 190244 112720 190256
rect 111852 190216 112720 190244
rect 111852 190204 111858 190216
rect 112714 190204 112720 190216
rect 112772 190244 112778 190256
rect 146846 190244 146852 190256
rect 112772 190216 146852 190244
rect 112772 190204 112778 190216
rect 146846 190204 146852 190216
rect 146904 190204 146910 190256
rect 169386 190204 169392 190256
rect 169444 190244 169450 190256
rect 194870 190244 194876 190256
rect 169444 190216 194876 190244
rect 169444 190204 169450 190216
rect 194870 190204 194876 190216
rect 194928 190204 194934 190256
rect 113174 190136 113180 190188
rect 113232 190176 113238 190188
rect 113726 190176 113732 190188
rect 113232 190148 113732 190176
rect 113232 190136 113238 190148
rect 113726 190136 113732 190148
rect 113784 190176 113790 190188
rect 146570 190176 146576 190188
rect 113784 190148 146576 190176
rect 113784 190136 113790 190148
rect 146570 190136 146576 190148
rect 146628 190136 146634 190188
rect 163498 190136 163504 190188
rect 163556 190176 163562 190188
rect 193674 190176 193680 190188
rect 163556 190148 193680 190176
rect 163556 190136 163562 190148
rect 193674 190136 193680 190148
rect 193732 190136 193738 190188
rect 111978 190068 111984 190120
rect 112036 190108 112042 190120
rect 145834 190108 145840 190120
rect 112036 190080 145840 190108
rect 112036 190068 112042 190080
rect 145834 190068 145840 190080
rect 145892 190068 145898 190120
rect 156690 190068 156696 190120
rect 156748 190108 156754 190120
rect 190914 190108 190920 190120
rect 156748 190080 190920 190108
rect 156748 190068 156754 190080
rect 190914 190068 190920 190080
rect 190972 190068 190978 190120
rect 111518 190000 111524 190052
rect 111576 190040 111582 190052
rect 136266 190040 136272 190052
rect 111576 190012 136272 190040
rect 111576 190000 111582 190012
rect 136266 190000 136272 190012
rect 136324 190000 136330 190052
rect 160646 190000 160652 190052
rect 160704 190040 160710 190052
rect 195146 190040 195152 190052
rect 160704 190012 195152 190040
rect 160704 190000 160710 190012
rect 195146 190000 195152 190012
rect 195204 190000 195210 190052
rect 109770 189932 109776 189984
rect 109828 189972 109834 189984
rect 133966 189972 133972 189984
rect 109828 189944 133972 189972
rect 109828 189932 109834 189944
rect 133966 189932 133972 189944
rect 134024 189932 134030 189984
rect 157518 189932 157524 189984
rect 157576 189972 157582 189984
rect 192478 189972 192484 189984
rect 157576 189944 192484 189972
rect 157576 189932 157582 189944
rect 192478 189932 192484 189944
rect 192536 189932 192542 189984
rect 119522 189864 119528 189916
rect 119580 189904 119586 189916
rect 150526 189904 150532 189916
rect 119580 189876 150532 189904
rect 119580 189864 119586 189876
rect 150526 189864 150532 189876
rect 150584 189864 150590 189916
rect 174170 189864 174176 189916
rect 174228 189904 174234 189916
rect 209222 189904 209228 189916
rect 174228 189876 209228 189904
rect 174228 189864 174234 189876
rect 209222 189864 209228 189876
rect 209280 189904 209286 189916
rect 260834 189904 260840 189916
rect 209280 189876 260840 189904
rect 209280 189864 209286 189876
rect 260834 189864 260840 189876
rect 260892 189864 260898 189916
rect 119706 189796 119712 189848
rect 119764 189836 119770 189848
rect 150986 189836 150992 189848
rect 119764 189808 150992 189836
rect 119764 189796 119770 189808
rect 150986 189796 150992 189808
rect 151044 189796 151050 189848
rect 157242 189796 157248 189848
rect 157300 189836 157306 189848
rect 192294 189836 192300 189848
rect 157300 189808 192300 189836
rect 157300 189796 157306 189808
rect 192294 189796 192300 189808
rect 192352 189796 192358 189848
rect 194870 189796 194876 189848
rect 194928 189836 194934 189848
rect 572254 189836 572260 189848
rect 194928 189808 572260 189836
rect 194928 189796 194934 189808
rect 572254 189796 572260 189808
rect 572312 189796 572318 189848
rect 107378 189728 107384 189780
rect 107436 189768 107442 189780
rect 139486 189768 139492 189780
rect 107436 189740 139492 189768
rect 107436 189728 107442 189740
rect 139486 189728 139492 189740
rect 139544 189728 139550 189780
rect 156414 189728 156420 189780
rect 156472 189768 156478 189780
rect 186130 189768 186136 189780
rect 156472 189740 186136 189768
rect 156472 189728 156478 189740
rect 186130 189728 186136 189740
rect 186188 189768 186194 189780
rect 579062 189768 579068 189780
rect 186188 189740 579068 189768
rect 186188 189728 186194 189740
rect 579062 189728 579068 189740
rect 579120 189728 579126 189780
rect 97350 189660 97356 189712
rect 97408 189700 97414 189712
rect 104894 189700 104900 189712
rect 97408 189672 104900 189700
rect 97408 189660 97414 189672
rect 104894 189660 104900 189672
rect 104952 189700 104958 189712
rect 149514 189700 149520 189712
rect 104952 189672 149520 189700
rect 104952 189660 104958 189672
rect 149514 189660 149520 189672
rect 149572 189660 149578 189712
rect 170306 189660 170312 189712
rect 170364 189700 170370 189712
rect 193214 189700 193220 189712
rect 170364 189672 193220 189700
rect 170364 189660 170370 189672
rect 193214 189660 193220 189672
rect 193272 189660 193278 189712
rect 111242 189592 111248 189644
rect 111300 189632 111306 189644
rect 142798 189632 142804 189644
rect 111300 189604 142804 189632
rect 111300 189592 111306 189604
rect 142798 189592 142804 189604
rect 142856 189592 142862 189644
rect 169294 189592 169300 189644
rect 169352 189632 169358 189644
rect 189074 189632 189080 189644
rect 169352 189604 189080 189632
rect 169352 189592 169358 189604
rect 189074 189592 189080 189604
rect 189132 189592 189138 189644
rect 170766 189524 170772 189576
rect 170824 189564 170830 189576
rect 189350 189564 189356 189576
rect 170824 189536 189356 189564
rect 170824 189524 170830 189536
rect 189350 189524 189356 189536
rect 189408 189524 189414 189576
rect 105814 189184 105820 189236
rect 105872 189224 105878 189236
rect 105872 189196 113174 189224
rect 105872 189184 105878 189196
rect 111978 189116 111984 189168
rect 112036 189156 112042 189168
rect 112438 189156 112444 189168
rect 112036 189128 112444 189156
rect 112036 189116 112042 189128
rect 112438 189116 112444 189128
rect 112496 189116 112502 189168
rect 113146 189156 113174 189196
rect 136634 189156 136640 189168
rect 113146 189128 136640 189156
rect 136634 189116 136640 189128
rect 136692 189116 136698 189168
rect 3418 189048 3424 189100
rect 3476 189088 3482 189100
rect 158622 189088 158628 189100
rect 3476 189060 158628 189088
rect 3476 189048 3482 189060
rect 158622 189048 158628 189060
rect 158680 189048 158686 189100
rect 206462 189048 206468 189100
rect 206520 189088 206526 189100
rect 579614 189088 579620 189100
rect 206520 189060 579620 189088
rect 206520 189048 206526 189060
rect 579614 189048 579620 189060
rect 579672 189048 579678 189100
rect 110414 188980 110420 189032
rect 110472 189020 110478 189032
rect 139854 189020 139860 189032
rect 110472 188992 139860 189020
rect 110472 188980 110478 188992
rect 139854 188980 139860 188992
rect 139912 188980 139918 189032
rect 144638 188980 144644 189032
rect 144696 189020 144702 189032
rect 570598 189020 570604 189032
rect 144696 188992 570604 189020
rect 144696 188980 144702 188992
rect 570598 188980 570604 188992
rect 570656 188980 570662 189032
rect 143442 188952 143448 188964
rect 142126 188924 143448 188952
rect 100018 188844 100024 188896
rect 100076 188884 100082 188896
rect 122926 188884 122932 188896
rect 100076 188856 122932 188884
rect 100076 188844 100082 188856
rect 122926 188844 122932 188856
rect 122984 188884 122990 188896
rect 123754 188884 123760 188896
rect 122984 188856 123760 188884
rect 122984 188844 122990 188856
rect 123754 188844 123760 188856
rect 123812 188844 123818 188896
rect 132126 188844 132132 188896
rect 132184 188884 132190 188896
rect 142126 188884 142154 188924
rect 143442 188912 143448 188924
rect 143500 188952 143506 188964
rect 568022 188952 568028 188964
rect 143500 188924 568028 188952
rect 143500 188912 143506 188924
rect 568022 188912 568028 188924
rect 568080 188912 568086 188964
rect 132184 188856 142154 188884
rect 132184 188844 132190 188856
rect 149698 188844 149704 188896
rect 149756 188884 149762 188896
rect 563790 188884 563796 188896
rect 149756 188856 563796 188884
rect 149756 188844 149762 188856
rect 563790 188844 563796 188856
rect 563848 188844 563854 188896
rect 94774 188776 94780 188828
rect 94832 188816 94838 188828
rect 126790 188816 126796 188828
rect 94832 188788 126796 188816
rect 94832 188776 94838 188788
rect 126790 188776 126796 188788
rect 126848 188776 126854 188828
rect 143442 188776 143448 188828
rect 143500 188816 143506 188828
rect 449158 188816 449164 188828
rect 143500 188788 449164 188816
rect 143500 188776 143506 188788
rect 449158 188776 449164 188788
rect 449216 188776 449222 188828
rect 94866 188708 94872 188760
rect 94924 188748 94930 188760
rect 110506 188748 110512 188760
rect 94924 188720 110512 188748
rect 94924 188708 94930 188720
rect 110506 188708 110512 188720
rect 110564 188708 110570 188760
rect 116854 188708 116860 188760
rect 116912 188748 116918 188760
rect 149698 188748 149704 188760
rect 116912 188720 149704 188748
rect 116912 188708 116918 188720
rect 149698 188708 149704 188720
rect 149756 188708 149762 188760
rect 150894 188708 150900 188760
rect 150952 188748 150958 188760
rect 269758 188748 269764 188760
rect 150952 188720 269764 188748
rect 150952 188708 150958 188720
rect 269758 188708 269764 188720
rect 269816 188708 269822 188760
rect 98730 188640 98736 188692
rect 98788 188680 98794 188692
rect 179414 188680 179420 188692
rect 98788 188652 179420 188680
rect 98788 188640 98794 188652
rect 179414 188640 179420 188652
rect 179472 188680 179478 188692
rect 205818 188680 205824 188692
rect 179472 188652 205824 188680
rect 179472 188640 179478 188652
rect 205818 188640 205824 188652
rect 205876 188640 205882 188692
rect 100294 188572 100300 188624
rect 100352 188612 100358 188624
rect 177206 188612 177212 188624
rect 100352 188584 177212 188612
rect 100352 188572 100358 188584
rect 177206 188572 177212 188584
rect 177264 188612 177270 188624
rect 207382 188612 207388 188624
rect 177264 188584 207388 188612
rect 177264 188572 177270 188584
rect 207382 188572 207388 188584
rect 207440 188572 207446 188624
rect 153102 188504 153108 188556
rect 153160 188544 153166 188556
rect 156874 188544 156880 188556
rect 153160 188516 156880 188544
rect 153160 188504 153166 188516
rect 156874 188504 156880 188516
rect 156932 188504 156938 188556
rect 171042 188504 171048 188556
rect 171100 188544 171106 188556
rect 206002 188544 206008 188556
rect 171100 188516 206008 188544
rect 171100 188504 171106 188516
rect 206002 188504 206008 188516
rect 206060 188544 206066 188556
rect 206462 188544 206468 188556
rect 206060 188516 206468 188544
rect 206060 188504 206066 188516
rect 206462 188504 206468 188516
rect 206520 188504 206526 188556
rect 95878 188436 95884 188488
rect 95936 188476 95942 188488
rect 154390 188476 154396 188488
rect 95936 188448 154396 188476
rect 95936 188436 95942 188448
rect 154390 188436 154396 188448
rect 154448 188436 154454 188488
rect 177758 188436 177764 188488
rect 177816 188476 177822 188488
rect 215846 188476 215852 188488
rect 177816 188448 215852 188476
rect 177816 188436 177822 188448
rect 215846 188436 215852 188448
rect 215904 188436 215910 188488
rect 89162 188368 89168 188420
rect 89220 188408 89226 188420
rect 153102 188408 153108 188420
rect 89220 188380 153108 188408
rect 89220 188368 89226 188380
rect 153102 188368 153108 188380
rect 153160 188368 153166 188420
rect 154316 188380 161474 188408
rect 53834 188300 53840 188352
rect 53892 188340 53898 188352
rect 107194 188340 107200 188352
rect 53892 188312 107200 188340
rect 53892 188300 53898 188312
rect 107194 188300 107200 188312
rect 107252 188300 107258 188352
rect 110506 188300 110512 188352
rect 110564 188340 110570 188352
rect 111426 188340 111432 188352
rect 110564 188312 111432 188340
rect 110564 188300 110570 188312
rect 111426 188300 111432 188312
rect 111484 188340 111490 188352
rect 145190 188340 145196 188352
rect 111484 188312 145196 188340
rect 111484 188300 111490 188312
rect 145190 188300 145196 188312
rect 145248 188300 145254 188352
rect 149514 188300 149520 188352
rect 149572 188340 149578 188352
rect 152734 188340 152740 188352
rect 149572 188312 152740 188340
rect 149572 188300 149578 188312
rect 152734 188300 152740 188312
rect 152792 188340 152798 188352
rect 154316 188340 154344 188380
rect 152792 188312 154344 188340
rect 161446 188340 161474 188380
rect 163222 188368 163228 188420
rect 163280 188408 163286 188420
rect 187050 188408 187056 188420
rect 163280 188380 187056 188408
rect 163280 188368 163286 188380
rect 187050 188368 187056 188380
rect 187108 188408 187114 188420
rect 241514 188408 241520 188420
rect 187108 188380 241520 188408
rect 187108 188368 187114 188380
rect 241514 188368 241520 188380
rect 241572 188368 241578 188420
rect 527174 188340 527180 188352
rect 161446 188312 527180 188340
rect 152792 188300 152798 188312
rect 527174 188300 527180 188312
rect 527232 188300 527238 188352
rect 123754 188232 123760 188284
rect 123812 188272 123818 188284
rect 155586 188272 155592 188284
rect 123812 188244 155592 188272
rect 123812 188232 123818 188244
rect 155586 188232 155592 188244
rect 155644 188232 155650 188284
rect 172882 188272 172888 188284
rect 161446 188244 172888 188272
rect 102778 188096 102784 188148
rect 102836 188136 102842 188148
rect 161446 188136 161474 188244
rect 172882 188232 172888 188244
rect 172940 188272 172946 188284
rect 203426 188272 203432 188284
rect 172940 188244 203432 188272
rect 172940 188232 172946 188244
rect 203426 188232 203432 188244
rect 203484 188232 203490 188284
rect 102836 188108 161474 188136
rect 102836 188096 102842 188108
rect 142798 187960 142804 188012
rect 142856 188000 142862 188012
rect 150894 188000 150900 188012
rect 142856 187972 150900 188000
rect 142856 187960 142862 187972
rect 150894 187960 150900 187972
rect 150952 187960 150958 188012
rect 105630 187756 105636 187808
rect 105688 187796 105694 187808
rect 110414 187796 110420 187808
rect 105688 187768 110420 187796
rect 105688 187756 105694 187768
rect 110414 187756 110420 187768
rect 110472 187756 110478 187808
rect 132034 187756 132040 187808
rect 132092 187796 132098 187808
rect 143442 187796 143448 187808
rect 132092 187768 143448 187796
rect 132092 187756 132098 187768
rect 143442 187756 143448 187768
rect 143500 187756 143506 187808
rect 154390 187756 154396 187808
rect 154448 187796 154454 187808
rect 155126 187796 155132 187808
rect 154448 187768 155132 187796
rect 154448 187756 154454 187768
rect 155126 187756 155132 187768
rect 155184 187756 155190 187808
rect 109586 187688 109592 187740
rect 109644 187728 109650 187740
rect 144638 187728 144644 187740
rect 109644 187700 144644 187728
rect 109644 187688 109650 187700
rect 144638 187688 144644 187700
rect 144696 187688 144702 187740
rect 91830 187620 91836 187672
rect 91888 187660 91894 187672
rect 171962 187660 171968 187672
rect 91888 187632 171968 187660
rect 91888 187620 91894 187632
rect 171962 187620 171968 187632
rect 172020 187660 172026 187672
rect 172238 187660 172244 187672
rect 172020 187632 172244 187660
rect 172020 187620 172026 187632
rect 172238 187620 172244 187632
rect 172296 187620 172302 187672
rect 199378 187620 199384 187672
rect 199436 187660 199442 187672
rect 200298 187660 200304 187672
rect 199436 187632 200304 187660
rect 199436 187620 199442 187632
rect 200298 187620 200304 187632
rect 200356 187660 200362 187672
rect 569218 187660 569224 187672
rect 200356 187632 569224 187660
rect 200356 187620 200362 187632
rect 569218 187620 569224 187632
rect 569276 187620 569282 187672
rect 84838 187552 84844 187604
rect 84896 187592 84902 187604
rect 84896 187564 142154 187592
rect 84896 187552 84902 187564
rect 107194 187484 107200 187536
rect 107252 187524 107258 187536
rect 136174 187524 136180 187536
rect 107252 187496 136180 187524
rect 107252 187484 107258 187496
rect 136174 187484 136180 187496
rect 136232 187484 136238 187536
rect 142126 187524 142154 187564
rect 166626 187552 166632 187604
rect 166684 187592 166690 187604
rect 201126 187592 201132 187604
rect 166684 187564 201132 187592
rect 166684 187552 166690 187564
rect 201126 187552 201132 187564
rect 201184 187552 201190 187604
rect 163590 187524 163596 187536
rect 142126 187496 163596 187524
rect 163590 187484 163596 187496
rect 163648 187524 163654 187536
rect 164142 187524 164148 187536
rect 163648 187496 164148 187524
rect 163648 187484 163654 187496
rect 164142 187484 164148 187496
rect 164200 187484 164206 187536
rect 168926 187484 168932 187536
rect 168984 187524 168990 187536
rect 201770 187524 201776 187536
rect 168984 187496 201776 187524
rect 168984 187484 168990 187496
rect 201770 187484 201776 187496
rect 201828 187484 201834 187536
rect 126238 187416 126244 187468
rect 126296 187456 126302 187468
rect 126790 187456 126796 187468
rect 126296 187428 126796 187456
rect 126296 187416 126302 187428
rect 126790 187416 126796 187428
rect 126848 187456 126854 187468
rect 151078 187456 151084 187468
rect 126848 187428 151084 187456
rect 126848 187416 126854 187428
rect 151078 187416 151084 187428
rect 151136 187416 151142 187468
rect 167454 187416 167460 187468
rect 167512 187456 167518 187468
rect 201678 187456 201684 187468
rect 167512 187428 201684 187456
rect 167512 187416 167518 187428
rect 201678 187416 201684 187428
rect 201736 187416 201742 187468
rect 115106 187348 115112 187400
rect 115164 187388 115170 187400
rect 147030 187388 147036 187400
rect 115164 187360 147036 187388
rect 115164 187348 115170 187360
rect 147030 187348 147036 187360
rect 147088 187348 147094 187400
rect 166074 187348 166080 187400
rect 166132 187388 166138 187400
rect 200574 187388 200580 187400
rect 166132 187360 200580 187388
rect 166132 187348 166138 187360
rect 200574 187348 200580 187360
rect 200632 187388 200638 187400
rect 201402 187388 201408 187400
rect 200632 187360 201408 187388
rect 200632 187348 200638 187360
rect 201402 187348 201408 187360
rect 201460 187348 201466 187400
rect 108942 187280 108948 187332
rect 109000 187320 109006 187332
rect 142338 187320 142344 187332
rect 109000 187292 142344 187320
rect 109000 187280 109006 187292
rect 142338 187280 142344 187292
rect 142396 187280 142402 187332
rect 163682 187280 163688 187332
rect 163740 187320 163746 187332
rect 197998 187320 198004 187332
rect 163740 187292 198004 187320
rect 163740 187280 163746 187292
rect 197998 187280 198004 187292
rect 198056 187280 198062 187332
rect 111610 187212 111616 187264
rect 111668 187252 111674 187264
rect 145098 187252 145104 187264
rect 111668 187224 145104 187252
rect 111668 187212 111674 187224
rect 145098 187212 145104 187224
rect 145156 187212 145162 187264
rect 158622 187212 158628 187264
rect 158680 187252 158686 187264
rect 193858 187252 193864 187264
rect 158680 187224 193864 187252
rect 158680 187212 158686 187224
rect 193858 187212 193864 187224
rect 193916 187212 193922 187264
rect 108574 187144 108580 187196
rect 108632 187184 108638 187196
rect 143350 187184 143356 187196
rect 108632 187156 143356 187184
rect 108632 187144 108638 187156
rect 143350 187144 143356 187156
rect 143408 187144 143414 187196
rect 165522 187144 165528 187196
rect 165580 187184 165586 187196
rect 203150 187184 203156 187196
rect 165580 187156 203156 187184
rect 165580 187144 165586 187156
rect 203150 187144 203156 187156
rect 203208 187144 203214 187196
rect 112622 187076 112628 187128
rect 112680 187116 112686 187128
rect 146754 187116 146760 187128
rect 112680 187088 146760 187116
rect 112680 187076 112686 187088
rect 146754 187076 146760 187088
rect 146812 187076 146818 187128
rect 173434 187076 173440 187128
rect 173492 187116 173498 187128
rect 211798 187116 211804 187128
rect 173492 187088 211804 187116
rect 173492 187076 173498 187088
rect 211798 187076 211804 187088
rect 211856 187076 211862 187128
rect 100294 187008 100300 187060
rect 100352 187048 100358 187060
rect 134978 187048 134984 187060
rect 100352 187020 134984 187048
rect 100352 187008 100358 187020
rect 134978 187008 134984 187020
rect 135036 187008 135042 187060
rect 135806 187008 135812 187060
rect 135864 187048 135870 187060
rect 136174 187048 136180 187060
rect 135864 187020 136180 187048
rect 135864 187008 135870 187020
rect 136174 187008 136180 187020
rect 136232 187008 136238 187060
rect 158346 187008 158352 187060
rect 158404 187048 158410 187060
rect 181990 187048 181996 187060
rect 158404 187020 181996 187048
rect 158404 187008 158410 187020
rect 181990 187008 181996 187020
rect 182048 187048 182054 187060
rect 278038 187048 278044 187060
rect 182048 187020 278044 187048
rect 182048 187008 182054 187020
rect 278038 187008 278044 187020
rect 278096 187008 278102 187060
rect 90542 186940 90548 186992
rect 90600 186980 90606 186992
rect 158622 186980 158628 186992
rect 90600 186952 158628 186980
rect 90600 186940 90606 186952
rect 158622 186940 158628 186952
rect 158680 186940 158686 186992
rect 162210 186940 162216 186992
rect 162268 186980 162274 186992
rect 196526 186980 196532 186992
rect 162268 186952 196532 186980
rect 162268 186940 162274 186952
rect 196526 186940 196532 186952
rect 196584 186940 196590 186992
rect 201402 186940 201408 186992
rect 201460 186980 201466 186992
rect 572070 186980 572076 186992
rect 201460 186952 572076 186980
rect 201460 186940 201466 186952
rect 572070 186940 572076 186952
rect 572128 186940 572134 186992
rect 164142 186872 164148 186924
rect 164200 186912 164206 186924
rect 176746 186912 176752 186924
rect 164200 186884 176752 186912
rect 164200 186872 164206 186884
rect 176746 186872 176752 186884
rect 176804 186872 176810 186924
rect 210234 186912 210240 186924
rect 180766 186884 210240 186912
rect 177666 186804 177672 186856
rect 177724 186844 177730 186856
rect 180766 186844 180794 186884
rect 210234 186872 210240 186884
rect 210292 186872 210298 186924
rect 177724 186816 180794 186844
rect 177724 186804 177730 186816
rect 130838 186328 130844 186380
rect 130896 186368 130902 186380
rect 144178 186368 144184 186380
rect 130896 186340 144184 186368
rect 130896 186328 130902 186340
rect 144178 186328 144184 186340
rect 144236 186368 144242 186380
rect 144822 186368 144828 186380
rect 144236 186340 144828 186368
rect 144236 186328 144242 186340
rect 144822 186328 144828 186340
rect 144880 186328 144886 186380
rect 158622 186328 158628 186380
rect 158680 186368 158686 186380
rect 160002 186368 160008 186380
rect 158680 186340 160008 186368
rect 158680 186328 158686 186340
rect 160002 186328 160008 186340
rect 160060 186328 160066 186380
rect 102870 186260 102876 186312
rect 102928 186300 102934 186312
rect 104342 186300 104348 186312
rect 102928 186272 104348 186300
rect 102928 186260 102934 186272
rect 104342 186260 104348 186272
rect 104400 186260 104406 186312
rect 112346 186260 112352 186312
rect 112404 186300 112410 186312
rect 145650 186300 145656 186312
rect 112404 186272 145656 186300
rect 112404 186260 112410 186272
rect 145650 186260 145656 186272
rect 145708 186300 145714 186312
rect 569402 186300 569408 186312
rect 145708 186272 569408 186300
rect 145708 186260 145714 186272
rect 569402 186260 569408 186272
rect 569460 186260 569466 186312
rect 138014 186192 138020 186244
rect 138072 186232 138078 186244
rect 558454 186232 558460 186244
rect 138072 186204 558460 186232
rect 138072 186192 138078 186204
rect 558454 186192 558460 186204
rect 558512 186192 558518 186244
rect 90358 186124 90364 186176
rect 90416 186164 90422 186176
rect 121546 186164 121552 186176
rect 90416 186136 121552 186164
rect 90416 186124 90422 186136
rect 121546 186124 121552 186136
rect 121604 186124 121610 186176
rect 144822 186124 144828 186176
rect 144880 186164 144886 186176
rect 511994 186164 512000 186176
rect 144880 186136 512000 186164
rect 144880 186124 144886 186136
rect 511994 186124 512000 186136
rect 512052 186124 512058 186176
rect 8294 186056 8300 186108
rect 8352 186096 8358 186108
rect 168742 186096 168748 186108
rect 8352 186068 168748 186096
rect 8352 186056 8358 186068
rect 168742 186056 168748 186068
rect 168800 186056 168806 186108
rect 97810 185988 97816 186040
rect 97868 186028 97874 186040
rect 189258 186028 189264 186040
rect 97868 186000 189264 186028
rect 97868 185988 97874 186000
rect 189258 185988 189264 186000
rect 189316 186028 189322 186040
rect 189316 186000 190454 186028
rect 189316 185988 189322 186000
rect 89254 185920 89260 185972
rect 89312 185960 89318 185972
rect 178402 185960 178408 185972
rect 89312 185932 178408 185960
rect 89312 185920 89318 185932
rect 178402 185920 178408 185932
rect 178460 185960 178466 185972
rect 190426 185960 190454 186000
rect 203334 185960 203340 185972
rect 178460 185932 180794 185960
rect 190426 185932 203340 185960
rect 178460 185920 178466 185932
rect 86402 185852 86408 185904
rect 86460 185892 86466 185904
rect 161750 185892 161756 185904
rect 86460 185864 161756 185892
rect 86460 185852 86466 185864
rect 161750 185852 161756 185864
rect 161808 185892 161814 185904
rect 162670 185892 162676 185904
rect 161808 185864 162676 185892
rect 161808 185852 161814 185864
rect 162670 185852 162676 185864
rect 162728 185852 162734 185904
rect 180766 185892 180794 185932
rect 203334 185920 203340 185932
rect 203392 185920 203398 185972
rect 211706 185892 211712 185904
rect 180766 185864 211712 185892
rect 211706 185852 211712 185864
rect 211764 185852 211770 185904
rect 93210 185784 93216 185836
rect 93268 185824 93274 185836
rect 164694 185824 164700 185836
rect 93268 185796 164700 185824
rect 93268 185784 93274 185796
rect 164694 185784 164700 185796
rect 164752 185824 164758 185836
rect 170398 185824 170404 185836
rect 164752 185796 170404 185824
rect 164752 185784 164758 185796
rect 170398 185784 170404 185796
rect 170456 185784 170462 185836
rect 173802 185784 173808 185836
rect 173860 185824 173866 185836
rect 207014 185824 207020 185836
rect 173860 185796 207020 185824
rect 173860 185784 173866 185796
rect 207014 185784 207020 185796
rect 207072 185784 207078 185836
rect 107654 185716 107660 185768
rect 107712 185756 107718 185768
rect 169202 185756 169208 185768
rect 107712 185728 169208 185756
rect 107712 185716 107718 185728
rect 169202 185716 169208 185728
rect 169260 185756 169266 185768
rect 211246 185756 211252 185768
rect 169260 185728 211252 185756
rect 169260 185716 169266 185728
rect 211246 185716 211252 185728
rect 211304 185716 211310 185768
rect 212442 185716 212448 185768
rect 212500 185756 212506 185768
rect 248414 185756 248420 185768
rect 212500 185728 248420 185756
rect 212500 185716 212506 185728
rect 248414 185716 248420 185728
rect 248472 185716 248478 185768
rect 104342 185648 104348 185700
rect 104400 185688 104406 185700
rect 138290 185688 138296 185700
rect 104400 185660 138296 185688
rect 104400 185648 104406 185660
rect 138290 185648 138296 185660
rect 138348 185648 138354 185700
rect 150710 185648 150716 185700
rect 150768 185688 150774 185700
rect 218422 185688 218428 185700
rect 150768 185660 218428 185688
rect 150768 185648 150774 185660
rect 218422 185648 218428 185660
rect 218480 185688 218486 185700
rect 306374 185688 306380 185700
rect 218480 185660 306380 185688
rect 218480 185648 218486 185660
rect 306374 185648 306380 185660
rect 306432 185648 306438 185700
rect 98822 185580 98828 185632
rect 98880 185620 98886 185632
rect 138014 185620 138020 185632
rect 98880 185592 138020 185620
rect 98880 185580 98886 185592
rect 138014 185580 138020 185592
rect 138072 185580 138078 185632
rect 147582 185580 147588 185632
rect 147640 185620 147646 185632
rect 215938 185620 215944 185632
rect 147640 185592 215944 185620
rect 147640 185580 147646 185592
rect 215938 185580 215944 185592
rect 215996 185620 216002 185632
rect 566734 185620 566740 185632
rect 215996 185592 566740 185620
rect 215996 185580 216002 185592
rect 566734 185580 566740 185592
rect 566792 185580 566798 185632
rect 106826 185512 106832 185564
rect 106884 185552 106890 185564
rect 108482 185552 108488 185564
rect 106884 185524 108488 185552
rect 106884 185512 106890 185524
rect 108482 185512 108488 185524
rect 108540 185552 108546 185564
rect 140406 185552 140412 185564
rect 108540 185524 140412 185552
rect 108540 185512 108546 185524
rect 140406 185512 140412 185524
rect 140464 185512 140470 185564
rect 160554 185512 160560 185564
rect 160612 185552 160618 185564
rect 211338 185552 211344 185564
rect 160612 185524 211344 185552
rect 160612 185512 160618 185524
rect 211338 185512 211344 185524
rect 211396 185552 211402 185564
rect 212442 185552 212448 185564
rect 211396 185524 212448 185552
rect 211396 185512 211402 185524
rect 212442 185512 212448 185524
rect 212500 185512 212506 185564
rect 121546 185444 121552 185496
rect 121604 185484 121610 185496
rect 121914 185484 121920 185496
rect 121604 185456 121920 185484
rect 121604 185444 121610 185456
rect 121914 185444 121920 185456
rect 121972 185484 121978 185496
rect 161474 185484 161480 185496
rect 121972 185456 161480 185484
rect 121972 185444 121978 185456
rect 161474 185444 161480 185456
rect 161532 185444 161538 185496
rect 3418 185104 3424 185156
rect 3476 185144 3482 185156
rect 7558 185144 7564 185156
rect 3476 185116 7564 185144
rect 3476 185104 3482 185116
rect 7558 185104 7564 185116
rect 7616 185104 7622 185156
rect 175642 184968 175648 185020
rect 175700 185008 175706 185020
rect 210418 185008 210424 185020
rect 175700 184980 210424 185008
rect 175700 184968 175706 184980
rect 210418 184968 210424 184980
rect 210476 184968 210482 185020
rect 168742 184900 168748 184952
rect 168800 184940 168806 184952
rect 210142 184940 210148 184952
rect 168800 184912 210148 184940
rect 168800 184900 168806 184912
rect 210142 184900 210148 184912
rect 210200 184900 210206 184952
rect 110322 184832 110328 184884
rect 110380 184872 110386 184884
rect 143810 184872 143816 184884
rect 110380 184844 143816 184872
rect 110380 184832 110386 184844
rect 143810 184832 143816 184844
rect 143868 184832 143874 184884
rect 144730 184832 144736 184884
rect 144788 184872 144794 184884
rect 581822 184872 581828 184884
rect 144788 184844 581828 184872
rect 144788 184832 144794 184844
rect 581822 184832 581828 184844
rect 581880 184832 581886 184884
rect 144822 184764 144828 184816
rect 144880 184804 144886 184816
rect 572346 184804 572352 184816
rect 144880 184776 572352 184804
rect 144880 184764 144886 184776
rect 572346 184764 572352 184776
rect 572404 184764 572410 184816
rect 98914 184696 98920 184748
rect 98972 184736 98978 184748
rect 167638 184736 167644 184748
rect 98972 184708 167644 184736
rect 98972 184696 98978 184708
rect 167638 184696 167644 184708
rect 167696 184736 167702 184748
rect 168190 184736 168196 184748
rect 167696 184708 168196 184736
rect 167696 184696 167702 184708
rect 168190 184696 168196 184708
rect 168248 184696 168254 184748
rect 173342 184696 173348 184748
rect 173400 184736 173406 184748
rect 204530 184736 204536 184748
rect 173400 184708 204536 184736
rect 173400 184696 173406 184708
rect 204530 184696 204536 184708
rect 204588 184696 204594 184748
rect 95970 184628 95976 184680
rect 96028 184668 96034 184680
rect 164602 184668 164608 184680
rect 96028 184640 164608 184668
rect 96028 184628 96034 184640
rect 164602 184628 164608 184640
rect 164660 184668 164666 184680
rect 165522 184668 165528 184680
rect 164660 184640 165528 184668
rect 164660 184628 164666 184640
rect 165522 184628 165528 184640
rect 165580 184628 165586 184680
rect 169938 184628 169944 184680
rect 169996 184668 170002 184680
rect 203886 184668 203892 184680
rect 169996 184640 203892 184668
rect 169996 184628 170002 184640
rect 203886 184628 203892 184640
rect 203944 184628 203950 184680
rect 101490 184560 101496 184612
rect 101548 184600 101554 184612
rect 168742 184600 168748 184612
rect 101548 184572 168748 184600
rect 101548 184560 101554 184572
rect 168742 184560 168748 184572
rect 168800 184560 168806 184612
rect 172238 184560 172244 184612
rect 172296 184600 172302 184612
rect 205726 184600 205732 184612
rect 172296 184572 205732 184600
rect 172296 184560 172302 184572
rect 205726 184560 205732 184572
rect 205784 184560 205790 184612
rect 99926 184492 99932 184544
rect 99984 184532 99990 184544
rect 158162 184532 158168 184544
rect 99984 184504 158168 184532
rect 99984 184492 99990 184504
rect 158162 184492 158168 184504
rect 158220 184492 158226 184544
rect 170030 184492 170036 184544
rect 170088 184532 170094 184544
rect 204622 184532 204628 184544
rect 170088 184504 204628 184532
rect 170088 184492 170094 184504
rect 204622 184492 204628 184504
rect 204680 184492 204686 184544
rect 121086 184424 121092 184476
rect 121144 184464 121150 184476
rect 154850 184464 154856 184476
rect 121144 184436 154856 184464
rect 121144 184424 121150 184436
rect 154850 184424 154856 184436
rect 154908 184424 154914 184476
rect 164878 184424 164884 184476
rect 164936 184464 164942 184476
rect 199010 184464 199016 184476
rect 164936 184436 199016 184464
rect 164936 184424 164942 184436
rect 199010 184424 199016 184436
rect 199068 184424 199074 184476
rect 105906 184356 105912 184408
rect 105964 184396 105970 184408
rect 139670 184396 139676 184408
rect 105964 184368 139676 184396
rect 105964 184356 105970 184368
rect 139670 184356 139676 184368
rect 139728 184356 139734 184408
rect 165430 184356 165436 184408
rect 165488 184396 165494 184408
rect 199286 184396 199292 184408
rect 165488 184368 199292 184396
rect 165488 184356 165494 184368
rect 199286 184356 199292 184368
rect 199344 184356 199350 184408
rect 110046 184288 110052 184340
rect 110104 184328 110110 184340
rect 143902 184328 143908 184340
rect 110104 184300 143908 184328
rect 110104 184288 110110 184300
rect 143902 184288 143908 184300
rect 143960 184288 143966 184340
rect 165522 184288 165528 184340
rect 165580 184328 165586 184340
rect 206094 184328 206100 184340
rect 165580 184300 206100 184328
rect 165580 184288 165586 184300
rect 206094 184288 206100 184300
rect 206152 184288 206158 184340
rect 109678 184220 109684 184272
rect 109736 184260 109742 184272
rect 143718 184260 143724 184272
rect 109736 184232 143724 184260
rect 109736 184220 109742 184232
rect 143718 184220 143724 184232
rect 143776 184260 143782 184272
rect 144822 184260 144828 184272
rect 143776 184232 144828 184260
rect 143776 184220 143782 184232
rect 144822 184220 144828 184232
rect 144880 184220 144886 184272
rect 159082 184220 159088 184272
rect 159140 184260 159146 184272
rect 181898 184260 181904 184272
rect 159140 184232 181904 184260
rect 159140 184220 159146 184232
rect 181898 184220 181904 184232
rect 181956 184260 181962 184272
rect 436094 184260 436100 184272
rect 181956 184232 436100 184260
rect 181956 184220 181962 184232
rect 436094 184220 436100 184232
rect 436152 184220 436158 184272
rect 109494 184152 109500 184204
rect 109552 184192 109558 184204
rect 144730 184192 144736 184204
rect 109552 184164 144736 184192
rect 109552 184152 109558 184164
rect 144730 184152 144736 184164
rect 144788 184152 144794 184204
rect 158254 184152 158260 184204
rect 158312 184192 158318 184204
rect 216950 184192 216956 184204
rect 158312 184164 216956 184192
rect 158312 184152 158318 184164
rect 216950 184152 216956 184164
rect 217008 184192 217014 184204
rect 563882 184192 563888 184204
rect 217008 184164 563888 184192
rect 217008 184152 217014 184164
rect 563882 184152 563888 184164
rect 563940 184152 563946 184204
rect 104342 184084 104348 184136
rect 104400 184124 104406 184136
rect 135898 184124 135904 184136
rect 104400 184096 135904 184124
rect 104400 184084 104406 184096
rect 135898 184084 135904 184096
rect 135956 184084 135962 184136
rect 160462 184084 160468 184136
rect 160520 184124 160526 184136
rect 190546 184124 190552 184136
rect 160520 184096 190552 184124
rect 160520 184084 160526 184096
rect 190546 184084 190552 184096
rect 190604 184084 190610 184136
rect 108758 184016 108764 184068
rect 108816 184056 108822 184068
rect 139578 184056 139584 184068
rect 108816 184028 139584 184056
rect 108816 184016 108822 184028
rect 139578 184016 139584 184028
rect 139636 184016 139642 184068
rect 176746 184016 176752 184068
rect 176804 184056 176810 184068
rect 204806 184056 204812 184068
rect 176804 184028 204812 184056
rect 176804 184016 176810 184028
rect 204806 184016 204812 184028
rect 204864 184016 204870 184068
rect 106090 183948 106096 184000
rect 106148 183988 106154 184000
rect 135530 183988 135536 184000
rect 106148 183960 135536 183988
rect 106148 183948 106154 183960
rect 135530 183948 135536 183960
rect 135588 183948 135594 184000
rect 168742 183948 168748 184000
rect 168800 183988 168806 184000
rect 188890 183988 188896 184000
rect 168800 183960 188896 183988
rect 168800 183948 168806 183960
rect 188890 183948 188896 183960
rect 188948 183948 188954 184000
rect 109954 183880 109960 183932
rect 110012 183920 110018 183932
rect 144546 183920 144552 183932
rect 110012 183892 144552 183920
rect 110012 183880 110018 183892
rect 144546 183880 144552 183892
rect 144604 183880 144610 183932
rect 80698 183472 80704 183524
rect 80756 183512 80762 183524
rect 178218 183512 178224 183524
rect 80756 183484 178224 183512
rect 80756 183472 80762 183484
rect 178218 183472 178224 183484
rect 178276 183512 178282 183524
rect 178402 183512 178408 183524
rect 178276 183484 178408 183512
rect 178276 183472 178282 183484
rect 178402 183472 178408 183484
rect 178460 183472 178466 183524
rect 101398 183404 101404 183456
rect 101456 183444 101462 183456
rect 178310 183444 178316 183456
rect 101456 183416 178316 183444
rect 101456 183404 101462 183416
rect 178310 183404 178316 183416
rect 178368 183404 178374 183456
rect 96154 183336 96160 183388
rect 96212 183376 96218 183388
rect 141142 183376 141148 183388
rect 96212 183348 141148 183376
rect 96212 183336 96218 183348
rect 141142 183336 141148 183348
rect 141200 183336 141206 183388
rect 156230 183336 156236 183388
rect 156288 183376 156294 183388
rect 202874 183376 202880 183388
rect 156288 183348 202880 183376
rect 156288 183336 156294 183348
rect 202874 183336 202880 183348
rect 202932 183376 202938 183388
rect 212994 183376 213000 183388
rect 202932 183348 213000 183376
rect 202932 183336 202938 183348
rect 212994 183336 213000 183348
rect 213052 183336 213058 183388
rect 178218 183268 178224 183320
rect 178276 183308 178282 183320
rect 212902 183308 212908 183320
rect 178276 183280 212908 183308
rect 178276 183268 178282 183280
rect 212902 183268 212908 183280
rect 212960 183268 212966 183320
rect 178310 183200 178316 183252
rect 178368 183240 178374 183252
rect 213086 183240 213092 183252
rect 178368 183212 213092 183240
rect 178368 183200 178374 183212
rect 213086 183200 213092 183212
rect 213144 183200 213150 183252
rect 165982 183132 165988 183184
rect 166040 183172 166046 183184
rect 207198 183172 207204 183184
rect 166040 183144 207204 183172
rect 166040 183132 166046 183144
rect 207198 183132 207204 183144
rect 207256 183132 207262 183184
rect 164510 183064 164516 183116
rect 164568 183104 164574 183116
rect 219618 183104 219624 183116
rect 164568 183076 219624 183104
rect 164568 183064 164574 183076
rect 219618 183064 219624 183076
rect 219676 183064 219682 183116
rect 159818 182996 159824 183048
rect 159876 183036 159882 183048
rect 219802 183036 219808 183048
rect 159876 183008 219808 183036
rect 159876 182996 159882 183008
rect 219802 182996 219808 183008
rect 219860 183036 219866 183048
rect 313274 183036 313280 183048
rect 219860 183008 313280 183036
rect 219860 182996 219866 183008
rect 313274 182996 313280 183008
rect 313332 182996 313338 183048
rect 156322 182928 156328 182980
rect 156380 182968 156386 182980
rect 216674 182968 216680 182980
rect 156380 182940 216680 182968
rect 156380 182928 156386 182940
rect 216674 182928 216680 182940
rect 216732 182968 216738 182980
rect 566826 182968 566832 182980
rect 216732 182940 566832 182968
rect 216732 182928 216738 182940
rect 566826 182928 566832 182940
rect 566884 182928 566890 182980
rect 158530 182860 158536 182912
rect 158588 182900 158594 182912
rect 215754 182900 215760 182912
rect 158588 182872 215760 182900
rect 158588 182860 158594 182872
rect 215754 182860 215760 182872
rect 215812 182900 215818 182912
rect 582374 182900 582380 182912
rect 215812 182872 582380 182900
rect 215812 182860 215818 182872
rect 582374 182860 582380 182872
rect 582432 182860 582438 182912
rect 86310 182792 86316 182844
rect 86368 182832 86374 182844
rect 125686 182832 125692 182844
rect 86368 182804 125692 182832
rect 86368 182792 86374 182804
rect 125686 182792 125692 182804
rect 125744 182832 125750 182844
rect 139210 182832 139216 182844
rect 125744 182804 139216 182832
rect 125744 182792 125750 182804
rect 139210 182792 139216 182804
rect 139268 182792 139274 182844
rect 153378 182792 153384 182844
rect 153436 182832 153442 182844
rect 214834 182832 214840 182844
rect 153436 182804 214840 182832
rect 153436 182792 153442 182804
rect 214834 182792 214840 182804
rect 214892 182832 214898 182844
rect 583018 182832 583024 182844
rect 214892 182804 583024 182832
rect 214892 182792 214898 182804
rect 583018 182792 583024 182804
rect 583076 182792 583082 182844
rect 218238 182452 218244 182504
rect 218296 182492 218302 182504
rect 218422 182492 218428 182504
rect 218296 182464 218428 182492
rect 218296 182452 218302 182464
rect 218422 182452 218428 182464
rect 218480 182452 218486 182504
rect 107102 182180 107108 182232
rect 107160 182220 107166 182232
rect 107160 182192 132494 182220
rect 107160 182180 107166 182192
rect 132466 182016 132494 182192
rect 187510 182180 187516 182232
rect 187568 182220 187574 182232
rect 191926 182220 191932 182232
rect 187568 182192 191932 182220
rect 187568 182180 187574 182192
rect 191926 182180 191932 182192
rect 191984 182220 191990 182232
rect 193122 182220 193128 182232
rect 191984 182192 193128 182220
rect 191984 182180 191990 182192
rect 193122 182180 193128 182192
rect 193180 182180 193186 182232
rect 143442 182112 143448 182164
rect 143500 182152 143506 182164
rect 150618 182152 150624 182164
rect 143500 182124 150624 182152
rect 143500 182112 143506 182124
rect 150618 182112 150624 182124
rect 150676 182152 150682 182164
rect 561214 182152 561220 182164
rect 150676 182124 561220 182152
rect 150676 182112 150682 182124
rect 561214 182112 561220 182124
rect 561272 182112 561278 182164
rect 162670 182044 162676 182096
rect 162728 182084 162734 182096
rect 189442 182084 189448 182096
rect 162728 182056 189448 182084
rect 162728 182044 162734 182056
rect 189442 182044 189448 182056
rect 189500 182044 189506 182096
rect 193122 182044 193128 182096
rect 193180 182084 193186 182096
rect 580166 182084 580172 182096
rect 193180 182056 580172 182084
rect 193180 182044 193186 182056
rect 580166 182044 580172 182056
rect 580224 182044 580230 182096
rect 142062 182016 142068 182028
rect 132466 181988 142068 182016
rect 142062 181976 142068 181988
rect 142120 182016 142126 182028
rect 213914 182016 213920 182028
rect 142120 181988 213920 182016
rect 142120 181976 142126 181988
rect 213914 181976 213920 181988
rect 213972 181976 213978 182028
rect 171226 181908 171232 181960
rect 171284 181948 171290 181960
rect 205910 181948 205916 181960
rect 171284 181920 205916 181948
rect 171284 181908 171290 181920
rect 205910 181908 205916 181920
rect 205968 181908 205974 181960
rect 176838 181840 176844 181892
rect 176896 181880 176902 181892
rect 211614 181880 211620 181892
rect 176896 181852 211620 181880
rect 176896 181840 176902 181852
rect 211614 181840 211620 181852
rect 211672 181840 211678 181892
rect 152918 181772 152924 181824
rect 152976 181812 152982 181824
rect 189258 181812 189264 181824
rect 152976 181784 189264 181812
rect 152976 181772 152982 181784
rect 189258 181772 189264 181784
rect 189316 181772 189322 181824
rect 105998 181704 106004 181756
rect 106056 181744 106062 181756
rect 137094 181744 137100 181756
rect 106056 181716 137100 181744
rect 106056 181704 106062 181716
rect 137094 181704 137100 181716
rect 137152 181704 137158 181756
rect 156138 181704 156144 181756
rect 156196 181744 156202 181756
rect 215662 181744 215668 181756
rect 156196 181716 215668 181744
rect 156196 181704 156202 181716
rect 215662 181704 215668 181716
rect 215720 181744 215726 181756
rect 233234 181744 233240 181756
rect 215720 181716 233240 181744
rect 215720 181704 215726 181716
rect 233234 181704 233240 181716
rect 233292 181704 233298 181756
rect 104250 181636 104256 181688
rect 104308 181676 104314 181688
rect 137922 181676 137928 181688
rect 104308 181648 137928 181676
rect 104308 181636 104314 181648
rect 137922 181636 137928 181648
rect 137980 181636 137986 181688
rect 159174 181636 159180 181688
rect 159232 181676 159238 181688
rect 180702 181676 180708 181688
rect 159232 181648 180708 181676
rect 159232 181636 159238 181648
rect 180702 181636 180708 181648
rect 180760 181676 180766 181688
rect 356054 181676 356060 181688
rect 180760 181648 356060 181676
rect 180760 181636 180766 181648
rect 356054 181636 356060 181648
rect 356112 181636 356118 181688
rect 103146 181568 103152 181620
rect 103204 181608 103210 181620
rect 137554 181608 137560 181620
rect 103204 181580 137560 181608
rect 103204 181568 103210 181580
rect 137554 181568 137560 181580
rect 137612 181568 137618 181620
rect 151998 181568 152004 181620
rect 152056 181608 152062 181620
rect 218514 181608 218520 181620
rect 152056 181580 218520 181608
rect 152056 181568 152062 181580
rect 218514 181568 218520 181580
rect 218572 181608 218578 181620
rect 562410 181608 562416 181620
rect 218572 181580 562416 181608
rect 218572 181568 218578 181580
rect 562410 181568 562416 181580
rect 562468 181568 562474 181620
rect 108390 181500 108396 181552
rect 108448 181540 108454 181552
rect 142430 181540 142436 181552
rect 108448 181512 142436 181540
rect 108448 181500 108454 181512
rect 142430 181500 142436 181512
rect 142488 181500 142494 181552
rect 149422 181500 149428 181552
rect 149480 181540 149486 181552
rect 217410 181540 217416 181552
rect 149480 181512 217416 181540
rect 149480 181500 149486 181512
rect 217410 181500 217416 181512
rect 217468 181540 217474 181552
rect 564066 181540 564072 181552
rect 217468 181512 564072 181540
rect 217468 181500 217474 181512
rect 564066 181500 564072 181512
rect 564124 181500 564130 181552
rect 94774 181432 94780 181484
rect 94832 181472 94838 181484
rect 117958 181472 117964 181484
rect 94832 181444 117964 181472
rect 94832 181432 94838 181444
rect 117958 181432 117964 181444
rect 118016 181432 118022 181484
rect 126882 181432 126888 181484
rect 126940 181472 126946 181484
rect 552750 181472 552756 181484
rect 126940 181444 552756 181472
rect 126940 181432 126946 181444
rect 552750 181432 552756 181444
rect 552808 181432 552814 181484
rect 174078 181364 174084 181416
rect 174136 181404 174142 181416
rect 208762 181404 208768 181416
rect 174136 181376 208768 181404
rect 174136 181364 174142 181376
rect 208762 181364 208768 181376
rect 208820 181364 208826 181416
rect 175458 181296 175464 181348
rect 175516 181336 175522 181348
rect 210326 181336 210332 181348
rect 175516 181308 210332 181336
rect 175516 181296 175522 181308
rect 210326 181296 210332 181308
rect 210384 181296 210390 181348
rect 3418 180820 3424 180872
rect 3476 180860 3482 180872
rect 94774 180860 94780 180872
rect 3476 180832 94780 180860
rect 3476 180820 3482 180832
rect 94774 180820 94780 180832
rect 94832 180820 94838 180872
rect 103054 180820 103060 180872
rect 103112 180860 103118 180872
rect 127802 180860 127808 180872
rect 103112 180832 127808 180860
rect 103112 180820 103118 180832
rect 127802 180820 127808 180832
rect 127860 180860 127866 180872
rect 127860 180832 128308 180860
rect 127860 180820 127866 180832
rect 128280 180792 128308 180832
rect 563974 180792 563980 180804
rect 128280 180764 563980 180792
rect 563974 180752 563980 180764
rect 564032 180752 564038 180804
rect 556798 180724 556804 180736
rect 132466 180696 556804 180724
rect 124030 180616 124036 180668
rect 124088 180656 124094 180668
rect 132466 180656 132494 180696
rect 556798 180684 556804 180696
rect 556856 180684 556862 180736
rect 124088 180628 132494 180656
rect 124088 180616 124094 180628
rect 136174 180616 136180 180668
rect 136232 180656 136238 180668
rect 558546 180656 558552 180668
rect 136232 180628 558552 180656
rect 136232 180616 136238 180628
rect 558546 180616 558552 180628
rect 558604 180616 558610 180668
rect 137002 180548 137008 180600
rect 137060 180588 137066 180600
rect 558362 180588 558368 180600
rect 137060 180560 558368 180588
rect 137060 180548 137066 180560
rect 558362 180548 558368 180560
rect 558420 180548 558426 180600
rect 120718 180480 120724 180532
rect 120776 180520 120782 180532
rect 455414 180520 455420 180532
rect 120776 180492 455420 180520
rect 120776 180480 120782 180492
rect 455414 180480 455420 180492
rect 455472 180480 455478 180532
rect 136910 180412 136916 180464
rect 136968 180452 136974 180464
rect 362954 180452 362960 180464
rect 136968 180424 362960 180452
rect 136968 180412 136974 180424
rect 362954 180412 362960 180424
rect 363012 180412 363018 180464
rect 120994 180276 121000 180328
rect 121052 180316 121058 180328
rect 136174 180316 136180 180328
rect 121052 180288 136180 180316
rect 121052 180276 121058 180288
rect 136174 180276 136180 180288
rect 136232 180276 136238 180328
rect 117958 180208 117964 180260
rect 118016 180248 118022 180260
rect 149330 180248 149336 180260
rect 118016 180220 149336 180248
rect 118016 180208 118022 180220
rect 149330 180208 149336 180220
rect 149388 180208 149394 180260
rect 102962 180140 102968 180192
rect 103020 180180 103026 180192
rect 137002 180180 137008 180192
rect 103020 180152 137008 180180
rect 103020 180140 103026 180152
rect 137002 180140 137008 180152
rect 137060 180140 137066 180192
rect 167362 180140 167368 180192
rect 167420 180180 167426 180192
rect 208854 180180 208860 180192
rect 167420 180152 208860 180180
rect 167420 180140 167426 180152
rect 208854 180140 208860 180152
rect 208912 180140 208918 180192
rect 102870 180072 102876 180124
rect 102928 180112 102934 180124
rect 136910 180112 136916 180124
rect 102928 180084 136916 180112
rect 102928 180072 102934 180084
rect 136910 180072 136916 180084
rect 136968 180072 136974 180124
rect 168650 180072 168656 180124
rect 168708 180112 168714 180124
rect 219710 180112 219716 180124
rect 168708 180084 219716 180112
rect 168708 180072 168714 180084
rect 219710 180072 219716 180084
rect 219768 180072 219774 180124
rect 127710 179324 127716 179376
rect 127768 179364 127774 179376
rect 581638 179364 581644 179376
rect 127768 179336 581644 179364
rect 127768 179324 127774 179336
rect 581638 179324 581644 179336
rect 581696 179324 581702 179376
rect 133782 179256 133788 179308
rect 133840 179296 133846 179308
rect 578970 179296 578976 179308
rect 133840 179268 578976 179296
rect 133840 179256 133846 179268
rect 578970 179256 578976 179268
rect 579028 179256 579034 179308
rect 138750 179188 138756 179240
rect 138808 179228 138814 179240
rect 558178 179228 558184 179240
rect 138808 179200 558184 179228
rect 138808 179188 138814 179200
rect 558178 179188 558184 179200
rect 558236 179188 558242 179240
rect 124766 179120 124772 179172
rect 124824 179160 124830 179172
rect 139026 179160 139032 179172
rect 124824 179132 139032 179160
rect 124824 179120 124830 179132
rect 139026 179120 139032 179132
rect 139084 179160 139090 179172
rect 405734 179160 405740 179172
rect 139084 179132 405740 179160
rect 139084 179120 139090 179132
rect 405734 179120 405740 179132
rect 405792 179120 405798 179172
rect 124030 179052 124036 179104
rect 124088 179092 124094 179104
rect 321554 179092 321560 179104
rect 124088 179064 321560 179092
rect 124088 179052 124094 179064
rect 321554 179052 321560 179064
rect 321612 179052 321618 179104
rect 170398 178848 170404 178900
rect 170456 178888 170462 178900
rect 203242 178888 203248 178900
rect 170456 178860 203248 178888
rect 170456 178848 170462 178860
rect 203242 178848 203248 178860
rect 203300 178848 203306 178900
rect 167638 178780 167644 178832
rect 167696 178820 167702 178832
rect 201862 178820 201868 178832
rect 167696 178792 201868 178820
rect 167696 178780 167702 178792
rect 201862 178780 201868 178792
rect 201920 178780 201926 178832
rect 105722 178712 105728 178764
rect 105780 178752 105786 178764
rect 132862 178752 132868 178764
rect 105780 178724 132868 178752
rect 105780 178712 105786 178724
rect 132862 178712 132868 178724
rect 132920 178752 132926 178764
rect 133782 178752 133788 178764
rect 132920 178724 133788 178752
rect 132920 178712 132926 178724
rect 133782 178712 133788 178724
rect 133840 178712 133846 178764
rect 161658 178712 161664 178764
rect 161716 178752 161722 178764
rect 210050 178752 210056 178764
rect 161716 178724 210056 178752
rect 161716 178712 161722 178724
rect 210050 178712 210056 178724
rect 210108 178752 210114 178764
rect 577774 178752 577780 178764
rect 210108 178724 577780 178752
rect 210108 178712 210114 178724
rect 577774 178712 577780 178724
rect 577832 178712 577838 178764
rect 105538 178644 105544 178696
rect 105596 178684 105602 178696
rect 138750 178684 138756 178696
rect 105596 178656 138756 178684
rect 105596 178644 105602 178656
rect 138750 178644 138756 178656
rect 138808 178644 138814 178696
rect 164418 178644 164424 178696
rect 164476 178684 164482 178696
rect 180610 178684 180616 178696
rect 164476 178656 180616 178684
rect 164476 178644 164482 178656
rect 180610 178644 180616 178656
rect 180668 178684 180674 178696
rect 560938 178684 560944 178696
rect 180668 178656 560944 178684
rect 180668 178644 180674 178656
rect 560938 178644 560944 178656
rect 560996 178644 561002 178696
rect 133782 177964 133788 178016
rect 133840 178004 133846 178016
rect 555418 178004 555424 178016
rect 133840 177976 555424 178004
rect 133840 177964 133846 177976
rect 555418 177964 555424 177976
rect 555476 177964 555482 178016
rect 131114 177896 131120 177948
rect 131172 177936 131178 177948
rect 132402 177936 132408 177948
rect 131172 177908 132408 177936
rect 131172 177896 131178 177908
rect 132402 177896 132408 177908
rect 132460 177936 132466 177948
rect 554038 177936 554044 177948
rect 132460 177908 554044 177936
rect 132460 177896 132466 177908
rect 554038 177896 554044 177908
rect 554096 177896 554102 177948
rect 191190 177828 191196 177880
rect 191248 177868 191254 177880
rect 580166 177868 580172 177880
rect 191248 177840 580172 177868
rect 191248 177828 191254 177840
rect 580166 177828 580172 177840
rect 580224 177828 580230 177880
rect 136542 177760 136548 177812
rect 136600 177800 136606 177812
rect 358814 177800 358820 177812
rect 136600 177772 358820 177800
rect 136600 177760 136606 177772
rect 358814 177760 358820 177772
rect 358872 177760 358878 177812
rect 101582 177420 101588 177472
rect 101640 177460 101646 177472
rect 131114 177460 131120 177472
rect 101640 177432 131120 177460
rect 101640 177420 101646 177432
rect 131114 177420 131120 177432
rect 131172 177420 131178 177472
rect 98914 177352 98920 177404
rect 98972 177392 98978 177404
rect 132770 177392 132776 177404
rect 98972 177364 132776 177392
rect 98972 177352 98978 177364
rect 132770 177352 132776 177364
rect 132828 177392 132834 177404
rect 133782 177392 133788 177404
rect 132828 177364 133788 177392
rect 132828 177352 132834 177364
rect 133782 177352 133788 177364
rect 133840 177352 133846 177404
rect 101490 177284 101496 177336
rect 101548 177324 101554 177336
rect 136542 177324 136548 177336
rect 101548 177296 136548 177324
rect 101548 177284 101554 177296
rect 136542 177284 136548 177296
rect 136600 177284 136606 177336
rect 100110 176672 100116 176724
rect 100168 176712 100174 176724
rect 122190 176712 122196 176724
rect 100168 176684 122196 176712
rect 100168 176672 100174 176684
rect 122190 176672 122196 176684
rect 122248 176712 122254 176724
rect 122248 176684 122834 176712
rect 122248 176672 122254 176684
rect 122806 176508 122834 176684
rect 136450 176604 136456 176656
rect 136508 176644 136514 176656
rect 552842 176644 552848 176656
rect 136508 176616 552848 176644
rect 136508 176604 136514 176616
rect 552842 176604 552848 176616
rect 552900 176604 552906 176656
rect 140774 176536 140780 176588
rect 140832 176576 140838 176588
rect 141050 176576 141056 176588
rect 140832 176548 141056 176576
rect 140832 176536 140838 176548
rect 141050 176536 141056 176548
rect 141108 176576 141114 176588
rect 555510 176576 555516 176588
rect 141108 176548 555516 176576
rect 141108 176536 141114 176548
rect 555510 176536 555516 176548
rect 555568 176536 555574 176588
rect 395338 176508 395344 176520
rect 122806 176480 395344 176508
rect 395338 176468 395344 176480
rect 395396 176468 395402 176520
rect 120902 175992 120908 176044
rect 120960 176032 120966 176044
rect 140774 176032 140780 176044
rect 120960 176004 140780 176032
rect 120960 175992 120966 176004
rect 140774 175992 140780 176004
rect 140832 175992 140838 176044
rect 101674 175924 101680 175976
rect 101732 175964 101738 175976
rect 136450 175964 136456 175976
rect 101732 175936 136456 175964
rect 101732 175924 101738 175936
rect 136450 175924 136456 175936
rect 136508 175924 136514 175976
rect 94866 173136 94872 173188
rect 94924 173176 94930 173188
rect 116486 173176 116492 173188
rect 94924 173148 116492 173176
rect 94924 173136 94930 173148
rect 116486 173136 116492 173148
rect 116544 173136 116550 173188
rect 185670 173136 185676 173188
rect 185728 173176 185734 173188
rect 580166 173176 580172 173188
rect 185728 173148 580172 173176
rect 185728 173136 185734 173148
rect 580166 173136 580172 173148
rect 580224 173136 580230 173188
rect 3418 172524 3424 172576
rect 3476 172564 3482 172576
rect 94682 172564 94688 172576
rect 3476 172536 94688 172564
rect 3476 172524 3482 172536
rect 94682 172524 94688 172536
rect 94740 172564 94746 172576
rect 94866 172564 94872 172576
rect 94740 172536 94872 172564
rect 94740 172524 94746 172536
rect 94866 172524 94872 172536
rect 94924 172524 94930 172576
rect 116486 171776 116492 171828
rect 116544 171816 116550 171828
rect 148778 171816 148784 171828
rect 116544 171788 148784 171816
rect 116544 171776 116550 171788
rect 148778 171776 148784 171788
rect 148836 171776 148842 171828
rect 110414 168988 110420 169040
rect 110472 169028 110478 169040
rect 111150 169028 111156 169040
rect 110472 169000 111156 169028
rect 110472 168988 110478 169000
rect 111150 168988 111156 169000
rect 111208 169028 111214 169040
rect 116394 169028 116400 169040
rect 111208 169000 116400 169028
rect 111208 168988 111214 169000
rect 116394 168988 116400 169000
rect 116452 168988 116458 169040
rect 3142 168376 3148 168428
rect 3200 168416 3206 168428
rect 110414 168416 110420 168428
rect 3200 168388 110420 168416
rect 3200 168376 3206 168388
rect 110414 168376 110420 168388
rect 110472 168376 110478 168428
rect 2774 165316 2780 165368
rect 2832 165356 2838 165368
rect 4798 165356 4804 165368
rect 2832 165328 4804 165356
rect 2832 165316 2838 165328
rect 4798 165316 4804 165328
rect 4856 165316 4862 165368
rect 188338 164228 188344 164280
rect 188396 164268 188402 164280
rect 580166 164268 580172 164280
rect 188396 164240 580172 164268
rect 188396 164228 188402 164240
rect 580166 164228 580172 164240
rect 580224 164228 580230 164280
rect 192570 162120 192576 162172
rect 192628 162160 192634 162172
rect 206186 162160 206192 162172
rect 192628 162132 206192 162160
rect 192628 162120 192634 162132
rect 206186 162120 206192 162132
rect 206244 162120 206250 162172
rect 206186 161440 206192 161492
rect 206244 161480 206250 161492
rect 580166 161480 580172 161492
rect 206244 161452 580172 161480
rect 206244 161440 206250 161452
rect 580166 161440 580172 161452
rect 580224 161440 580230 161492
rect 3510 161372 3516 161424
rect 3568 161412 3574 161424
rect 171134 161412 171140 161424
rect 3568 161384 171140 161412
rect 3568 161372 3574 161384
rect 171134 161372 171140 161384
rect 171192 161412 171198 161424
rect 172238 161412 172244 161424
rect 171192 161384 172244 161412
rect 171192 161372 171198 161384
rect 172238 161372 172244 161384
rect 172296 161372 172302 161424
rect 172238 160692 172244 160744
rect 172296 160732 172302 160744
rect 191926 160732 191932 160744
rect 172296 160704 191932 160732
rect 172296 160692 172302 160704
rect 191926 160692 191932 160704
rect 191984 160692 191990 160744
rect 3510 155932 3516 155984
rect 3568 155972 3574 155984
rect 116946 155972 116952 155984
rect 3568 155944 116952 155972
rect 3568 155932 3574 155944
rect 116946 155932 116952 155944
rect 117004 155972 117010 155984
rect 117004 155944 117268 155972
rect 117004 155932 117010 155944
rect 117240 155904 117268 155944
rect 127618 155904 127624 155916
rect 117240 155876 127624 155904
rect 127618 155864 127624 155876
rect 127676 155864 127682 155916
rect 163130 153824 163136 153876
rect 163188 153864 163194 153876
rect 198090 153864 198096 153876
rect 163188 153836 198096 153864
rect 163188 153824 163194 153836
rect 198090 153824 198096 153836
rect 198148 153824 198154 153876
rect 198090 153212 198096 153264
rect 198148 153252 198154 153264
rect 579614 153252 579620 153264
rect 198148 153224 579620 153252
rect 198148 153212 198154 153224
rect 579614 153212 579620 153224
rect 579672 153212 579678 153264
rect 113542 153144 113548 153196
rect 113600 153184 113606 153196
rect 117774 153184 117780 153196
rect 113600 153156 117780 153184
rect 113600 153144 113606 153156
rect 117774 153144 117780 153156
rect 117832 153144 117838 153196
rect 3510 151784 3516 151836
rect 3568 151824 3574 151836
rect 113542 151824 113548 151836
rect 3568 151796 113548 151824
rect 3568 151784 3574 151796
rect 113542 151784 113548 151796
rect 113600 151784 113606 151836
rect 99926 151240 99932 151292
rect 99984 151280 99990 151292
rect 132678 151280 132684 151292
rect 99984 151252 132684 151280
rect 99984 151240 99990 151252
rect 132678 151240 132684 151252
rect 132736 151240 132742 151292
rect 175458 151240 175464 151292
rect 175516 151280 175522 151292
rect 210602 151280 210608 151292
rect 175516 151252 210608 151280
rect 175516 151240 175522 151252
rect 210602 151240 210608 151252
rect 210660 151240 210666 151292
rect 100018 151172 100024 151224
rect 100076 151212 100082 151224
rect 134334 151212 134340 151224
rect 100076 151184 134340 151212
rect 100076 151172 100082 151184
rect 134334 151172 134340 151184
rect 134392 151172 134398 151224
rect 165890 151172 165896 151224
rect 165948 151212 165954 151224
rect 217502 151212 217508 151224
rect 165948 151184 217508 151212
rect 165948 151172 165954 151184
rect 217502 151172 217508 151184
rect 217560 151172 217566 151224
rect 98638 151104 98644 151156
rect 98696 151144 98702 151156
rect 132586 151144 132592 151156
rect 98696 151116 132592 151144
rect 98696 151104 98702 151116
rect 132586 151104 132592 151116
rect 132644 151104 132650 151156
rect 154758 151104 154764 151156
rect 154816 151144 154822 151156
rect 214558 151144 214564 151156
rect 154816 151116 214564 151144
rect 154816 151104 154822 151116
rect 214558 151104 214564 151116
rect 214616 151104 214622 151156
rect 99834 151036 99840 151088
rect 99892 151076 99898 151088
rect 134058 151076 134064 151088
rect 99892 151048 134064 151076
rect 99892 151036 99898 151048
rect 134058 151036 134064 151048
rect 134116 151036 134122 151088
rect 156046 151036 156052 151088
rect 156104 151076 156110 151088
rect 216030 151076 216036 151088
rect 156104 151048 216036 151076
rect 156104 151036 156110 151048
rect 216030 151036 216036 151048
rect 216088 151036 216094 151088
rect 214650 149676 214656 149728
rect 214708 149716 214714 149728
rect 580166 149716 580172 149728
rect 214708 149688 580172 149716
rect 214708 149676 214714 149688
rect 580166 149676 580172 149688
rect 580224 149676 580230 149728
rect 3418 148996 3424 149048
rect 3476 149036 3482 149048
rect 160370 149036 160376 149048
rect 3476 149008 160376 149036
rect 3476 148996 3482 149008
rect 160370 148996 160376 149008
rect 160428 149036 160434 149048
rect 160428 149008 161474 149036
rect 160428 148996 160434 149008
rect 106918 148928 106924 148980
rect 106976 148968 106982 148980
rect 132310 148968 132316 148980
rect 106976 148940 132316 148968
rect 106976 148928 106982 148940
rect 132310 148928 132316 148940
rect 132368 148928 132374 148980
rect 161446 148968 161474 149008
rect 173986 148996 173992 149048
rect 174044 149036 174050 149048
rect 207658 149036 207664 149048
rect 174044 149008 207664 149036
rect 174044 148996 174050 149008
rect 207658 148996 207664 149008
rect 207716 148996 207722 149048
rect 194778 148968 194784 148980
rect 161446 148940 194784 148968
rect 194778 148928 194784 148940
rect 194836 148928 194842 148980
rect 106826 148860 106832 148912
rect 106884 148900 106890 148912
rect 132218 148900 132224 148912
rect 106884 148872 132224 148900
rect 106884 148860 106890 148872
rect 132218 148860 132224 148872
rect 132276 148860 132282 148912
rect 165246 148860 165252 148912
rect 165304 148900 165310 148912
rect 199654 148900 199660 148912
rect 165304 148872 199660 148900
rect 165304 148860 165310 148872
rect 199654 148860 199660 148872
rect 199712 148860 199718 148912
rect 104066 148792 104072 148844
rect 104124 148832 104130 148844
rect 133230 148832 133236 148844
rect 104124 148804 133236 148832
rect 104124 148792 104130 148804
rect 133230 148792 133236 148804
rect 133288 148792 133294 148844
rect 163038 148792 163044 148844
rect 163096 148832 163102 148844
rect 198274 148832 198280 148844
rect 163096 148804 198280 148832
rect 163096 148792 163102 148804
rect 198274 148792 198280 148804
rect 198332 148792 198338 148844
rect 110690 148724 110696 148776
rect 110748 148764 110754 148776
rect 144454 148764 144460 148776
rect 110748 148736 144460 148764
rect 110748 148724 110754 148736
rect 144454 148724 144460 148736
rect 144512 148724 144518 148776
rect 167270 148724 167276 148776
rect 167328 148764 167334 148776
rect 201954 148764 201960 148776
rect 167328 148736 201960 148764
rect 167328 148724 167334 148736
rect 201954 148724 201960 148736
rect 202012 148724 202018 148776
rect 101214 148656 101220 148708
rect 101272 148696 101278 148708
rect 134242 148696 134248 148708
rect 101272 148668 134248 148696
rect 101272 148656 101278 148668
rect 134242 148656 134248 148668
rect 134300 148656 134306 148708
rect 161566 148656 161572 148708
rect 161624 148696 161630 148708
rect 196894 148696 196900 148708
rect 161624 148668 196900 148696
rect 161624 148656 161630 148668
rect 196894 148656 196900 148668
rect 196952 148656 196958 148708
rect 98730 148588 98736 148640
rect 98788 148628 98794 148640
rect 132954 148628 132960 148640
rect 98788 148600 132960 148628
rect 98788 148588 98794 148600
rect 132954 148588 132960 148600
rect 133012 148588 133018 148640
rect 168098 148588 168104 148640
rect 168156 148628 168162 148640
rect 202046 148628 202052 148640
rect 168156 148600 202052 148628
rect 168156 148588 168162 148600
rect 202046 148588 202052 148600
rect 202104 148588 202110 148640
rect 108298 148520 108304 148572
rect 108356 148560 108362 148572
rect 142614 148560 142620 148572
rect 108356 148532 142620 148560
rect 108356 148520 108362 148532
rect 142614 148520 142620 148532
rect 142672 148520 142678 148572
rect 168558 148520 168564 148572
rect 168616 148560 168622 148572
rect 203610 148560 203616 148572
rect 168616 148532 203616 148560
rect 168616 148520 168622 148532
rect 203610 148520 203616 148532
rect 203668 148520 203674 148572
rect 101398 148452 101404 148504
rect 101456 148492 101462 148504
rect 135714 148492 135720 148504
rect 101456 148464 135720 148492
rect 101456 148452 101462 148464
rect 135714 148452 135720 148464
rect 135772 148452 135778 148504
rect 169846 148452 169852 148504
rect 169904 148492 169910 148504
rect 204990 148492 204996 148504
rect 169904 148464 204996 148492
rect 169904 148452 169910 148464
rect 204990 148452 204996 148464
rect 205048 148452 205054 148504
rect 107010 148384 107016 148436
rect 107068 148424 107074 148436
rect 143994 148424 144000 148436
rect 107068 148396 144000 148424
rect 107068 148384 107074 148396
rect 143994 148384 144000 148396
rect 144052 148384 144058 148436
rect 175366 148384 175372 148436
rect 175424 148424 175430 148436
rect 211982 148424 211988 148436
rect 175424 148396 211988 148424
rect 175424 148384 175430 148396
rect 211982 148384 211988 148396
rect 212040 148384 212046 148436
rect 97902 148316 97908 148368
rect 97960 148356 97966 148368
rect 131758 148356 131764 148368
rect 97960 148328 131764 148356
rect 97960 148316 97966 148328
rect 131758 148316 131764 148328
rect 131816 148316 131822 148368
rect 174630 148316 174636 148368
rect 174688 148356 174694 148368
rect 211890 148356 211896 148368
rect 174688 148328 211896 148356
rect 174688 148316 174694 148328
rect 211890 148316 211896 148328
rect 211948 148316 211954 148368
rect 120810 148248 120816 148300
rect 120868 148288 120874 148300
rect 141694 148288 141700 148300
rect 120868 148260 141700 148288
rect 120868 148248 120874 148260
rect 141694 148248 141700 148260
rect 141752 148248 141758 148300
rect 167178 148248 167184 148300
rect 167236 148288 167242 148300
rect 200666 148288 200672 148300
rect 167236 148260 200672 148288
rect 167236 148248 167242 148260
rect 200666 148248 200672 148260
rect 200724 148248 200730 148300
rect 110782 148180 110788 148232
rect 110840 148220 110846 148232
rect 130746 148220 130752 148232
rect 110840 148192 130752 148220
rect 110840 148180 110846 148192
rect 130746 148180 130752 148192
rect 130804 148180 130810 148232
rect 172330 148180 172336 148232
rect 172388 148220 172394 148232
rect 202138 148220 202144 148232
rect 172388 148192 202144 148220
rect 172388 148180 172394 148192
rect 202138 148180 202144 148192
rect 202196 148180 202202 148232
rect 114830 148112 114836 148164
rect 114888 148152 114894 148164
rect 130654 148152 130660 148164
rect 114888 148124 130660 148152
rect 114888 148112 114894 148124
rect 130654 148112 130660 148124
rect 130712 148112 130718 148164
rect 180242 148112 180248 148164
rect 180300 148152 180306 148164
rect 192754 148152 192760 148164
rect 180300 148124 192760 148152
rect 180300 148112 180306 148124
rect 192754 148112 192760 148124
rect 192812 148112 192818 148164
rect 171870 147296 171876 147348
rect 171928 147336 171934 147348
rect 189810 147336 189816 147348
rect 171928 147308 189816 147336
rect 171928 147296 171934 147308
rect 189810 147296 189816 147308
rect 189868 147296 189874 147348
rect 176194 147228 176200 147280
rect 176252 147268 176258 147280
rect 196066 147268 196072 147280
rect 176252 147240 196072 147268
rect 176252 147228 176258 147240
rect 196066 147228 196072 147240
rect 196124 147228 196130 147280
rect 168006 147160 168012 147212
rect 168064 147200 168070 147212
rect 194042 147200 194048 147212
rect 168064 147172 194048 147200
rect 168064 147160 168070 147172
rect 194042 147160 194048 147172
rect 194100 147160 194106 147212
rect 165798 147092 165804 147144
rect 165856 147132 165862 147144
rect 201402 147132 201408 147144
rect 165856 147104 201408 147132
rect 165856 147092 165862 147104
rect 201402 147092 201408 147104
rect 201460 147092 201466 147144
rect 112162 147024 112168 147076
rect 112220 147064 112226 147076
rect 140314 147064 140320 147076
rect 112220 147036 140320 147064
rect 112220 147024 112226 147036
rect 140314 147024 140320 147036
rect 140372 147024 140378 147076
rect 165706 147024 165712 147076
rect 165764 147064 165770 147076
rect 206370 147064 206376 147076
rect 165764 147036 206376 147064
rect 165764 147024 165770 147036
rect 206370 147024 206376 147036
rect 206428 147024 206434 147076
rect 101306 146956 101312 147008
rect 101364 146996 101370 147008
rect 135622 146996 135628 147008
rect 101364 146968 135628 146996
rect 101364 146956 101370 146968
rect 135622 146956 135628 146968
rect 135680 146956 135686 147008
rect 168374 146956 168380 147008
rect 168432 146996 168438 147008
rect 210510 146996 210516 147008
rect 168432 146968 210516 146996
rect 168432 146956 168438 146968
rect 210510 146956 210516 146968
rect 210568 146956 210574 147008
rect 102686 146888 102692 146940
rect 102744 146928 102750 146940
rect 137462 146928 137468 146940
rect 102744 146900 137468 146928
rect 102744 146888 102750 146900
rect 137462 146888 137468 146900
rect 137520 146928 137526 146940
rect 580166 146928 580172 146940
rect 137520 146900 580172 146928
rect 137520 146888 137526 146900
rect 580166 146888 580172 146900
rect 580224 146888 580230 146940
rect 183278 146820 183284 146872
rect 183336 146860 183342 146872
rect 183462 146860 183468 146872
rect 183336 146832 183468 146860
rect 183336 146820 183342 146832
rect 183462 146820 183468 146832
rect 183520 146820 183526 146872
rect 200942 146276 200948 146328
rect 201000 146316 201006 146328
rect 201402 146316 201408 146328
rect 201000 146288 201408 146316
rect 201000 146276 201006 146288
rect 201402 146276 201408 146288
rect 201460 146316 201466 146328
rect 580442 146316 580448 146328
rect 201460 146288 580448 146316
rect 201460 146276 201466 146288
rect 580442 146276 580448 146288
rect 580500 146276 580506 146328
rect 116670 146208 116676 146260
rect 116728 146248 116734 146260
rect 129366 146248 129372 146260
rect 116728 146220 129372 146248
rect 116728 146208 116734 146220
rect 129366 146208 129372 146220
rect 129424 146208 129430 146260
rect 179874 146208 179880 146260
rect 179932 146248 179938 146260
rect 197906 146248 197912 146260
rect 179932 146220 197912 146248
rect 179932 146208 179938 146220
rect 197906 146208 197912 146220
rect 197964 146208 197970 146260
rect 115198 146140 115204 146192
rect 115256 146180 115262 146192
rect 127066 146180 127072 146192
rect 115256 146152 127072 146180
rect 115256 146140 115262 146152
rect 127066 146140 127072 146152
rect 127124 146140 127130 146192
rect 177574 146140 177580 146192
rect 177632 146180 177638 146192
rect 199746 146180 199752 146192
rect 177632 146152 199752 146180
rect 177632 146140 177638 146152
rect 199746 146140 199752 146152
rect 199804 146140 199810 146192
rect 113450 146072 113456 146124
rect 113508 146112 113514 146124
rect 130378 146112 130384 146124
rect 113508 146084 130384 146112
rect 113508 146072 113514 146084
rect 130378 146072 130384 146084
rect 130436 146072 130442 146124
rect 173986 146072 173992 146124
rect 174044 146112 174050 146124
rect 199102 146112 199108 146124
rect 174044 146084 199108 146112
rect 174044 146072 174050 146084
rect 199102 146072 199108 146084
rect 199160 146072 199166 146124
rect 112530 146004 112536 146056
rect 112588 146044 112594 146056
rect 131758 146044 131764 146056
rect 112588 146016 131764 146044
rect 112588 146004 112594 146016
rect 131758 146004 131764 146016
rect 131816 146004 131822 146056
rect 172606 146004 172612 146056
rect 172664 146044 172670 146056
rect 197814 146044 197820 146056
rect 172664 146016 197820 146044
rect 172664 146004 172670 146016
rect 197814 146004 197820 146016
rect 197872 146004 197878 146056
rect 114186 145936 114192 145988
rect 114244 145976 114250 145988
rect 134242 145976 134248 145988
rect 114244 145948 134248 145976
rect 114244 145936 114250 145948
rect 134242 145936 134248 145948
rect 134300 145936 134306 145988
rect 162946 145936 162952 145988
rect 163004 145976 163010 145988
rect 188338 145976 188344 145988
rect 163004 145948 188344 145976
rect 163004 145936 163010 145948
rect 188338 145936 188344 145948
rect 188396 145936 188402 145988
rect 111702 145868 111708 145920
rect 111760 145908 111766 145920
rect 135254 145908 135260 145920
rect 111760 145880 135260 145908
rect 111760 145868 111766 145880
rect 135254 145868 135260 145880
rect 135312 145868 135318 145920
rect 169846 145868 169852 145920
rect 169904 145908 169910 145920
rect 198734 145908 198740 145920
rect 169904 145880 198740 145908
rect 169904 145868 169910 145880
rect 198734 145868 198740 145880
rect 198792 145868 198798 145920
rect 112898 145800 112904 145852
rect 112956 145840 112962 145852
rect 144086 145840 144092 145852
rect 112956 145812 144092 145840
rect 112956 145800 112962 145812
rect 144086 145800 144092 145812
rect 144144 145800 144150 145852
rect 167362 145800 167368 145852
rect 167420 145840 167426 145852
rect 198918 145840 198924 145852
rect 167420 145812 198924 145840
rect 167420 145800 167426 145812
rect 198918 145800 198924 145812
rect 198976 145800 198982 145852
rect 119246 145732 119252 145784
rect 119304 145772 119310 145784
rect 153746 145772 153752 145784
rect 119304 145744 153752 145772
rect 119304 145732 119310 145744
rect 153746 145732 153752 145744
rect 153804 145732 153810 145784
rect 160370 145732 160376 145784
rect 160428 145772 160434 145784
rect 193582 145772 193588 145784
rect 160428 145744 193588 145772
rect 160428 145732 160434 145744
rect 193582 145732 193588 145744
rect 193640 145732 193646 145784
rect 118142 145664 118148 145716
rect 118200 145704 118206 145716
rect 151906 145704 151912 145716
rect 118200 145676 151912 145704
rect 118200 145664 118206 145676
rect 151906 145664 151912 145676
rect 151964 145664 151970 145716
rect 164326 145664 164332 145716
rect 164384 145704 164390 145716
rect 197630 145704 197636 145716
rect 164384 145676 197636 145704
rect 164384 145664 164390 145676
rect 197630 145664 197636 145676
rect 197688 145664 197694 145716
rect 119614 145596 119620 145648
rect 119672 145636 119678 145648
rect 154482 145636 154488 145648
rect 119672 145608 154488 145636
rect 119672 145596 119678 145608
rect 154482 145596 154488 145608
rect 154540 145596 154546 145648
rect 162394 145596 162400 145648
rect 162452 145636 162458 145648
rect 195238 145636 195244 145648
rect 162452 145608 195244 145636
rect 162452 145596 162458 145608
rect 195238 145596 195244 145608
rect 195296 145596 195302 145648
rect 117866 145528 117872 145580
rect 117924 145568 117930 145580
rect 152366 145568 152372 145580
rect 117924 145540 152372 145568
rect 117924 145528 117930 145540
rect 152366 145528 152372 145540
rect 152424 145528 152430 145580
rect 162486 145528 162492 145580
rect 162544 145568 162550 145580
rect 196802 145568 196808 145580
rect 162544 145540 196808 145568
rect 162544 145528 162550 145540
rect 196802 145528 196808 145540
rect 196860 145528 196866 145580
rect 112898 145460 112904 145512
rect 112956 145500 112962 145512
rect 124214 145500 124220 145512
rect 112956 145472 124220 145500
rect 112956 145460 112962 145472
rect 124214 145460 124220 145472
rect 124272 145460 124278 145512
rect 177298 145460 177304 145512
rect 177356 145500 177362 145512
rect 192386 145500 192392 145512
rect 177356 145472 192392 145500
rect 177356 145460 177362 145472
rect 192386 145460 192392 145472
rect 192444 145460 192450 145512
rect 116210 145392 116216 145444
rect 116268 145432 116274 145444
rect 122926 145432 122932 145444
rect 116268 145404 122932 145432
rect 116268 145392 116274 145404
rect 122926 145392 122932 145404
rect 122984 145392 122990 145444
rect 181438 145392 181444 145444
rect 181496 145432 181502 145444
rect 196250 145432 196256 145444
rect 181496 145404 196256 145432
rect 181496 145392 181502 145404
rect 196250 145392 196256 145404
rect 196308 145392 196314 145444
rect 113818 145324 113824 145376
rect 113876 145364 113882 145376
rect 125226 145364 125232 145376
rect 113876 145336 125232 145364
rect 113876 145324 113882 145336
rect 125226 145324 125232 145336
rect 125284 145324 125290 145376
rect 184934 145324 184940 145376
rect 184992 145364 184998 145376
rect 196434 145364 196440 145376
rect 184992 145336 196440 145364
rect 184992 145324 184998 145336
rect 196434 145324 196440 145336
rect 196492 145324 196498 145376
rect 120626 145256 120632 145308
rect 120684 145296 120690 145308
rect 121362 145296 121368 145308
rect 120684 145268 121368 145296
rect 120684 145256 120690 145268
rect 121362 145256 121368 145268
rect 121420 145256 121426 145308
rect 188246 144984 188252 145036
rect 188304 145024 188310 145036
rect 188890 145024 188896 145036
rect 188304 144996 188896 145024
rect 188304 144984 188310 144996
rect 188890 144984 188896 144996
rect 188948 144984 188954 145036
rect 3418 144916 3424 144968
rect 3476 144956 3482 144968
rect 119062 144956 119068 144968
rect 3476 144928 119068 144956
rect 3476 144916 3482 144928
rect 119062 144916 119068 144928
rect 119120 144956 119126 144968
rect 119246 144956 119252 144968
rect 119120 144928 119252 144956
rect 119120 144916 119126 144928
rect 119246 144916 119252 144928
rect 119304 144916 119310 144968
rect 3510 144848 3516 144900
rect 3568 144888 3574 144900
rect 113910 144888 113916 144900
rect 3568 144860 113916 144888
rect 3568 144848 3574 144860
rect 113910 144848 113916 144860
rect 113968 144888 113974 144900
rect 114186 144888 114192 144900
rect 113968 144860 114192 144888
rect 113968 144848 113974 144860
rect 114186 144848 114192 144860
rect 114244 144848 114250 144900
rect 121822 144848 121828 144900
rect 121880 144888 121886 144900
rect 138658 144888 138664 144900
rect 121880 144860 138664 144888
rect 121880 144848 121886 144860
rect 138658 144848 138664 144860
rect 138716 144848 138722 144900
rect 176654 144848 176660 144900
rect 176712 144888 176718 144900
rect 196342 144888 196348 144900
rect 176712 144860 196348 144888
rect 176712 144848 176718 144860
rect 196342 144848 196348 144860
rect 196400 144848 196406 144900
rect 197538 144848 197544 144900
rect 197596 144888 197602 144900
rect 197722 144888 197728 144900
rect 197596 144860 197728 144888
rect 197596 144848 197602 144860
rect 197722 144848 197728 144860
rect 197780 144888 197786 144900
rect 580258 144888 580264 144900
rect 197780 144860 580264 144888
rect 197780 144848 197786 144860
rect 580258 144848 580264 144860
rect 580316 144848 580322 144900
rect 110966 144780 110972 144832
rect 111024 144820 111030 144832
rect 130562 144820 130568 144832
rect 111024 144792 130568 144820
rect 111024 144780 111030 144792
rect 130562 144780 130568 144792
rect 130620 144780 130626 144832
rect 175274 144780 175280 144832
rect 175332 144820 175338 144832
rect 199562 144820 199568 144832
rect 175332 144792 199568 144820
rect 175332 144780 175338 144792
rect 199562 144780 199568 144792
rect 199620 144780 199626 144832
rect 114462 144712 114468 144764
rect 114520 144752 114526 144764
rect 140130 144752 140136 144764
rect 114520 144724 140136 144752
rect 114520 144712 114526 144724
rect 140130 144712 140136 144724
rect 140188 144712 140194 144764
rect 166902 144712 166908 144764
rect 166960 144752 166966 144764
rect 196250 144752 196256 144764
rect 166960 144724 196256 144752
rect 166960 144712 166966 144724
rect 196250 144712 196256 144724
rect 196308 144712 196314 144764
rect 114278 144644 114284 144696
rect 114336 144684 114342 144696
rect 141786 144684 141792 144696
rect 114336 144656 141792 144684
rect 114336 144644 114342 144656
rect 141786 144644 141792 144656
rect 141844 144644 141850 144696
rect 157334 144644 157340 144696
rect 157392 144684 157398 144696
rect 189534 144684 189540 144696
rect 157392 144656 189540 144684
rect 157392 144644 157398 144656
rect 189534 144644 189540 144656
rect 189592 144644 189598 144696
rect 115566 144576 115572 144628
rect 115624 144616 115630 144628
rect 142890 144616 142896 144628
rect 115624 144588 142896 144616
rect 115624 144576 115630 144588
rect 142890 144576 142896 144588
rect 142948 144576 142954 144628
rect 158162 144576 158168 144628
rect 158220 144616 158226 144628
rect 190822 144616 190828 144628
rect 158220 144588 190828 144616
rect 158220 144576 158226 144588
rect 190822 144576 190828 144588
rect 190880 144576 190886 144628
rect 117682 144508 117688 144560
rect 117740 144548 117746 144560
rect 149882 144548 149888 144560
rect 117740 144520 149888 144548
rect 117740 144508 117746 144520
rect 149882 144508 149888 144520
rect 149940 144508 149946 144560
rect 160278 144508 160284 144560
rect 160336 144548 160342 144560
rect 195514 144548 195520 144560
rect 160336 144520 195520 144548
rect 160336 144508 160342 144520
rect 195514 144508 195520 144520
rect 195572 144508 195578 144560
rect 116394 144440 116400 144492
rect 116452 144480 116458 144492
rect 148410 144480 148416 144492
rect 116452 144452 148416 144480
rect 116452 144440 116458 144452
rect 148410 144440 148416 144452
rect 148468 144440 148474 144492
rect 160186 144440 160192 144492
rect 160244 144480 160250 144492
rect 194870 144480 194876 144492
rect 160244 144452 194876 144480
rect 160244 144440 160250 144452
rect 194870 144440 194876 144452
rect 194928 144440 194934 144492
rect 114738 144372 114744 144424
rect 114796 144412 114802 144424
rect 148870 144412 148876 144424
rect 114796 144384 148876 144412
rect 114796 144372 114802 144384
rect 148870 144372 148876 144384
rect 148928 144372 148934 144424
rect 161290 144372 161296 144424
rect 161348 144412 161354 144424
rect 195606 144412 195612 144424
rect 161348 144384 195612 144412
rect 161348 144372 161354 144384
rect 195606 144372 195612 144384
rect 195664 144372 195670 144424
rect 111334 144304 111340 144356
rect 111392 144344 111398 144356
rect 145190 144344 145196 144356
rect 111392 144316 145196 144344
rect 111392 144304 111398 144316
rect 145190 144304 145196 144316
rect 145248 144304 145254 144356
rect 158070 144304 158076 144356
rect 158128 144344 158134 144356
rect 194226 144344 194232 144356
rect 158128 144316 194232 144344
rect 158128 144304 158134 144316
rect 194226 144304 194232 144316
rect 194284 144304 194290 144356
rect 111702 144236 111708 144288
rect 111760 144276 111766 144288
rect 146294 144276 146300 144288
rect 111760 144248 146300 144276
rect 111760 144236 111766 144248
rect 146294 144236 146300 144248
rect 146352 144236 146358 144288
rect 155862 144236 155868 144288
rect 155920 144276 155926 144288
rect 191834 144276 191840 144288
rect 155920 144248 191840 144276
rect 155920 144236 155926 144248
rect 191834 144236 191840 144248
rect 191892 144236 191898 144288
rect 112990 144168 112996 144220
rect 113048 144208 113054 144220
rect 137922 144208 137928 144220
rect 113048 144180 137928 144208
rect 113048 144168 113054 144180
rect 137922 144168 137928 144180
rect 137980 144208 137986 144220
rect 188154 144208 188160 144220
rect 137980 144180 188160 144208
rect 137980 144168 137986 144180
rect 188154 144168 188160 144180
rect 188212 144168 188218 144220
rect 196250 144168 196256 144220
rect 196308 144208 196314 144220
rect 197078 144208 197084 144220
rect 196308 144180 197084 144208
rect 196308 144168 196314 144180
rect 197078 144168 197084 144180
rect 197136 144208 197142 144220
rect 207566 144208 207572 144220
rect 197136 144180 207572 144208
rect 197136 144168 197142 144180
rect 207566 144168 207572 144180
rect 207624 144168 207630 144220
rect 114186 144100 114192 144152
rect 114244 144140 114250 144152
rect 126974 144140 126980 144152
rect 114244 144112 126980 144140
rect 114244 144100 114250 144112
rect 126974 144100 126980 144112
rect 127032 144100 127038 144152
rect 177482 144100 177488 144152
rect 177540 144140 177546 144152
rect 198182 144140 198188 144152
rect 177540 144112 198188 144140
rect 177540 144100 177546 144112
rect 198182 144100 198188 144112
rect 198240 144100 198246 144152
rect 187602 144032 187608 144084
rect 187660 144072 187666 144084
rect 197538 144072 197544 144084
rect 187660 144044 197544 144072
rect 187660 144032 187666 144044
rect 197538 144032 197544 144044
rect 197596 144032 197602 144084
rect 121546 143664 121552 143676
rect 115906 143636 121552 143664
rect 97810 143556 97816 143608
rect 97868 143596 97874 143608
rect 97868 143568 110460 143596
rect 97868 143556 97874 143568
rect 110432 143528 110460 143568
rect 111058 143528 111064 143540
rect 110432 143500 111064 143528
rect 111058 143488 111064 143500
rect 111116 143528 111122 143540
rect 115906 143528 115934 143636
rect 121546 143624 121552 143636
rect 121604 143624 121610 143676
rect 191098 143624 191104 143676
rect 191156 143664 191162 143676
rect 534074 143664 534080 143676
rect 191156 143636 534080 143664
rect 191156 143624 191162 143636
rect 534074 143624 534080 143636
rect 534132 143624 534138 143676
rect 118418 143556 118424 143608
rect 118476 143596 118482 143608
rect 123662 143596 123668 143608
rect 118476 143568 123668 143596
rect 118476 143556 118482 143568
rect 123662 143556 123668 143568
rect 123720 143596 123726 143608
rect 492674 143596 492680 143608
rect 123720 143568 492680 143596
rect 123720 143556 123726 143568
rect 492674 143556 492680 143568
rect 492732 143556 492738 143608
rect 111116 143500 115934 143528
rect 121104 143500 121316 143528
rect 111116 143488 111122 143500
rect 115474 143420 115480 143472
rect 115532 143460 115538 143472
rect 121104 143460 121132 143500
rect 115532 143432 121132 143460
rect 121288 143460 121316 143500
rect 121454 143488 121460 143540
rect 121512 143528 121518 143540
rect 122190 143528 122196 143540
rect 121512 143500 122196 143528
rect 121512 143488 121518 143500
rect 122190 143488 122196 143500
rect 122248 143488 122254 143540
rect 122282 143488 122288 143540
rect 122340 143528 122346 143540
rect 127618 143528 127624 143540
rect 122340 143500 127624 143528
rect 122340 143488 122346 143500
rect 127618 143488 127624 143500
rect 127676 143488 127682 143540
rect 127728 143500 128354 143528
rect 127728 143460 127756 143500
rect 121288 143432 127756 143460
rect 128326 143460 128354 143500
rect 172514 143488 172520 143540
rect 172572 143528 172578 143540
rect 173710 143528 173716 143540
rect 172572 143500 173716 143528
rect 172572 143488 172578 143500
rect 173710 143488 173716 143500
rect 173768 143488 173774 143540
rect 133506 143460 133512 143472
rect 128326 143432 133512 143460
rect 115532 143420 115538 143432
rect 133506 143420 133512 143432
rect 133564 143420 133570 143472
rect 115198 143352 115204 143404
rect 115256 143392 115262 143404
rect 119890 143392 119896 143404
rect 115256 143364 119896 143392
rect 115256 143352 115262 143364
rect 119890 143352 119896 143364
rect 119948 143392 119954 143404
rect 119948 143364 121132 143392
rect 119948 143352 119954 143364
rect 97994 143216 98000 143268
rect 98052 143256 98058 143268
rect 98052 143228 115520 143256
rect 98052 143216 98058 143228
rect 97258 142944 97264 142996
rect 97316 142984 97322 142996
rect 115198 142984 115204 142996
rect 97316 142956 115204 142984
rect 97316 142944 97322 142956
rect 115198 142944 115204 142956
rect 115256 142944 115262 142996
rect 82814 142808 82820 142860
rect 82872 142848 82878 142860
rect 115492 142848 115520 143228
rect 116302 143216 116308 143268
rect 116360 143256 116366 143268
rect 116670 143256 116676 143268
rect 116360 143228 116676 143256
rect 116360 143216 116366 143228
rect 116670 143216 116676 143228
rect 116728 143256 116734 143268
rect 121104 143256 121132 143364
rect 121546 143352 121552 143404
rect 121604 143392 121610 143404
rect 127710 143392 127716 143404
rect 121604 143364 127716 143392
rect 121604 143352 121610 143364
rect 127710 143352 127716 143364
rect 127768 143352 127774 143404
rect 127802 143352 127808 143404
rect 127860 143392 127866 143404
rect 138566 143392 138572 143404
rect 127860 143364 138572 143392
rect 127860 143352 127866 143364
rect 138566 143352 138572 143364
rect 138624 143352 138630 143404
rect 179322 143352 179328 143404
rect 179380 143392 179386 143404
rect 187602 143392 187608 143404
rect 179380 143364 187608 143392
rect 179380 143352 179386 143364
rect 187602 143352 187608 143364
rect 187660 143352 187666 143404
rect 121362 143284 121368 143336
rect 121420 143324 121426 143336
rect 139394 143324 139400 143336
rect 121420 143296 139400 143324
rect 121420 143284 121426 143296
rect 139394 143284 139400 143296
rect 139452 143284 139458 143336
rect 181346 143284 181352 143336
rect 181404 143324 181410 143336
rect 192018 143324 192024 143336
rect 181404 143296 192024 143324
rect 181404 143284 181410 143296
rect 192018 143284 192024 143296
rect 192076 143284 192082 143336
rect 122282 143256 122288 143268
rect 116728 143228 120580 143256
rect 121104 143228 122288 143256
rect 116728 143216 116734 143228
rect 115658 143148 115664 143200
rect 115716 143188 115722 143200
rect 120442 143188 120448 143200
rect 115716 143160 120448 143188
rect 115716 143148 115722 143160
rect 120442 143148 120448 143160
rect 120500 143148 120506 143200
rect 120552 143188 120580 143228
rect 122282 143216 122288 143228
rect 122340 143216 122346 143268
rect 126974 143216 126980 143268
rect 127032 143256 127038 143268
rect 147674 143256 147680 143268
rect 127032 143228 147680 143256
rect 127032 143216 127038 143228
rect 147674 143216 147680 143228
rect 147732 143216 147738 143268
rect 177206 143216 177212 143268
rect 177264 143256 177270 143268
rect 195054 143256 195060 143268
rect 177264 143228 195060 143256
rect 177264 143216 177270 143228
rect 195054 143216 195060 143228
rect 195112 143216 195118 143268
rect 140958 143188 140964 143200
rect 120552 143160 140964 143188
rect 140958 143148 140964 143160
rect 141016 143148 141022 143200
rect 175182 143148 175188 143200
rect 175240 143188 175246 143200
rect 197630 143188 197636 143200
rect 175240 143160 197636 143188
rect 175240 143148 175246 143160
rect 197630 143148 197636 143160
rect 197688 143188 197694 143200
rect 197688 143160 200114 143188
rect 197688 143148 197694 143160
rect 118510 143080 118516 143132
rect 118568 143120 118574 143132
rect 145926 143120 145932 143132
rect 118568 143092 118694 143120
rect 118568 143080 118574 143092
rect 118666 143052 118694 143092
rect 120552 143092 145932 143120
rect 120552 143052 120580 143092
rect 145926 143080 145932 143092
rect 145984 143080 145990 143132
rect 163866 143080 163872 143132
rect 163924 143120 163930 143132
rect 193490 143120 193496 143132
rect 163924 143092 193496 143120
rect 163924 143080 163930 143092
rect 193490 143080 193496 143092
rect 193548 143080 193554 143132
rect 118666 143024 120580 143052
rect 120626 143012 120632 143064
rect 120684 143052 120690 143064
rect 143534 143052 143540 143064
rect 120684 143024 143540 143052
rect 120684 143012 120690 143024
rect 143534 143012 143540 143024
rect 143592 143012 143598 143064
rect 162302 143012 162308 143064
rect 162360 143052 162366 143064
rect 194962 143052 194968 143064
rect 162360 143024 194968 143052
rect 162360 143012 162366 143024
rect 194962 143012 194968 143024
rect 195020 143012 195026 143064
rect 116578 142944 116584 142996
rect 116636 142984 116642 142996
rect 119890 142984 119896 142996
rect 116636 142956 119896 142984
rect 116636 142944 116642 142956
rect 119890 142944 119896 142956
rect 119948 142944 119954 142996
rect 119982 142944 119988 142996
rect 120040 142984 120046 142996
rect 150894 142984 150900 142996
rect 120040 142956 150900 142984
rect 120040 142944 120046 142956
rect 150894 142944 150900 142956
rect 150952 142944 150958 142996
rect 155678 142944 155684 142996
rect 155736 142984 155742 142996
rect 157334 142984 157340 142996
rect 155736 142956 157340 142984
rect 155736 142944 155742 142956
rect 157334 142944 157340 142956
rect 157392 142944 157398 142996
rect 159818 142944 159824 142996
rect 159876 142984 159882 142996
rect 193766 142984 193772 142996
rect 159876 142956 193772 142984
rect 159876 142944 159882 142956
rect 193766 142944 193772 142956
rect 193824 142944 193830 142996
rect 200086 142984 200114 143160
rect 270494 142984 270500 142996
rect 200086 142956 270500 142984
rect 270494 142944 270500 142956
rect 270552 142944 270558 142996
rect 116762 142876 116768 142928
rect 116820 142916 116826 142928
rect 149238 142916 149244 142928
rect 116820 142888 149244 142916
rect 116820 142876 116826 142888
rect 149238 142876 149244 142888
rect 149296 142876 149302 142928
rect 168926 142876 168932 142928
rect 168984 142916 168990 142928
rect 192202 142916 192208 142928
rect 168984 142888 192208 142916
rect 168984 142876 168990 142888
rect 192202 142876 192208 142888
rect 192260 142876 192266 142928
rect 192386 142876 192392 142928
rect 192444 142916 192450 142928
rect 580258 142916 580264 142928
rect 192444 142888 580264 142916
rect 192444 142876 192450 142888
rect 580258 142876 580264 142888
rect 580316 142876 580322 142928
rect 119798 142848 119804 142860
rect 82872 142820 103514 142848
rect 115492 142820 119804 142848
rect 82872 142808 82878 142820
rect 103486 142780 103514 142820
rect 119798 142808 119804 142820
rect 119856 142808 119862 142860
rect 119890 142808 119896 142860
rect 119948 142848 119954 142860
rect 120074 142848 120080 142860
rect 119948 142820 120080 142848
rect 119948 142808 119954 142820
rect 120074 142808 120080 142820
rect 120132 142848 120138 142860
rect 121362 142848 121368 142860
rect 120132 142820 121368 142848
rect 120132 142808 120138 142820
rect 121362 142808 121368 142820
rect 121420 142808 121426 142860
rect 122282 142808 122288 142860
rect 122340 142848 122346 142860
rect 153378 142848 153384 142860
rect 122340 142820 153384 142848
rect 122340 142808 122346 142820
rect 153378 142808 153384 142820
rect 153436 142808 153442 142860
rect 166442 142808 166448 142860
rect 166500 142848 166506 142860
rect 169754 142848 169760 142860
rect 166500 142820 169760 142848
rect 166500 142808 166506 142820
rect 169754 142808 169760 142820
rect 169812 142808 169818 142860
rect 171042 142808 171048 142860
rect 171100 142848 171106 142860
rect 191098 142848 191104 142860
rect 171100 142820 191104 142848
rect 171100 142808 171106 142820
rect 191098 142808 191104 142820
rect 191156 142808 191162 142860
rect 192110 142808 192116 142860
rect 192168 142848 192174 142860
rect 580718 142848 580724 142860
rect 192168 142820 580724 142848
rect 192168 142808 192174 142820
rect 580718 142808 580724 142820
rect 580776 142808 580782 142860
rect 116670 142780 116676 142792
rect 103486 142752 116676 142780
rect 116670 142740 116676 142752
rect 116728 142740 116734 142792
rect 118234 142740 118240 142792
rect 118292 142780 118298 142792
rect 131114 142780 131120 142792
rect 118292 142752 131120 142780
rect 118292 142740 118298 142752
rect 131114 142740 131120 142752
rect 131172 142740 131178 142792
rect 173710 142740 173716 142792
rect 173768 142780 173774 142792
rect 179690 142780 179696 142792
rect 173768 142752 179696 142780
rect 173768 142740 173774 142752
rect 179690 142740 179696 142752
rect 179748 142740 179754 142792
rect 117130 142672 117136 142724
rect 117188 142712 117194 142724
rect 128538 142712 128544 142724
rect 117188 142684 128544 142712
rect 117188 142672 117194 142684
rect 128538 142672 128544 142684
rect 128596 142672 128602 142724
rect 176378 142672 176384 142724
rect 176436 142712 176442 142724
rect 178586 142712 178592 142724
rect 176436 142684 178592 142712
rect 176436 142672 176442 142684
rect 178586 142672 178592 142684
rect 178644 142672 178650 142724
rect 115750 142604 115756 142656
rect 115808 142644 115814 142656
rect 126054 142644 126060 142656
rect 115808 142616 126060 142644
rect 115808 142604 115814 142616
rect 126054 142604 126060 142616
rect 126112 142604 126118 142656
rect 131114 142604 131120 142656
rect 131172 142644 131178 142656
rect 426434 142644 426440 142656
rect 131172 142616 426440 142644
rect 131172 142604 131178 142616
rect 426434 142604 426440 142616
rect 426492 142604 426498 142656
rect 119798 142536 119804 142588
rect 119856 142576 119862 142588
rect 122282 142576 122288 142588
rect 119856 142548 122288 142576
rect 119856 142536 119862 142548
rect 122282 142536 122288 142548
rect 122340 142536 122346 142588
rect 154482 142536 154488 142588
rect 154540 142576 154546 142588
rect 514754 142576 514760 142588
rect 154540 142548 514760 142576
rect 154540 142536 154546 142548
rect 514754 142536 514760 142548
rect 514812 142536 514818 142588
rect 173710 142468 173716 142520
rect 173768 142508 173774 142520
rect 179414 142508 179420 142520
rect 173768 142480 179420 142508
rect 173768 142468 173774 142480
rect 179414 142468 179420 142480
rect 179472 142468 179478 142520
rect 179690 142468 179696 142520
rect 179748 142508 179754 142520
rect 207842 142508 207848 142520
rect 179748 142480 207848 142508
rect 179748 142468 179754 142480
rect 207842 142468 207848 142480
rect 207900 142468 207906 142520
rect 142890 142400 142896 142452
rect 142948 142440 142954 142452
rect 188982 142440 188988 142452
rect 142948 142412 188988 142440
rect 142948 142400 142954 142412
rect 188982 142400 188988 142412
rect 189040 142400 189046 142452
rect 59354 142332 59360 142384
rect 59412 142372 59418 142384
rect 177206 142372 177212 142384
rect 59412 142344 177212 142372
rect 59412 142332 59418 142344
rect 177206 142332 177212 142344
rect 177264 142332 177270 142384
rect 187602 142332 187608 142384
rect 187660 142372 187666 142384
rect 220814 142372 220820 142384
rect 187660 142344 220820 142372
rect 187660 142332 187666 142344
rect 220814 142332 220820 142344
rect 220872 142332 220878 142384
rect 152366 142264 152372 142316
rect 152424 142304 152430 142316
rect 365714 142304 365720 142316
rect 152424 142276 365720 142304
rect 152424 142264 152430 142276
rect 365714 142264 365720 142276
rect 365772 142264 365778 142316
rect 161382 142128 161388 142180
rect 161440 142168 161446 142180
rect 161440 142140 169064 142168
rect 161440 142128 161446 142140
rect 115906 142072 119844 142100
rect 114278 141992 114284 142044
rect 114336 142032 114342 142044
rect 115906 142032 115934 142072
rect 114336 142004 115934 142032
rect 119816 142032 119844 142072
rect 119890 142060 119896 142112
rect 119948 142100 119954 142112
rect 151446 142100 151452 142112
rect 119948 142072 151452 142100
rect 119948 142060 119954 142072
rect 151446 142060 151452 142072
rect 151504 142060 151510 142112
rect 169036 142100 169064 142140
rect 193306 142100 193312 142112
rect 169036 142072 193312 142100
rect 193306 142060 193312 142072
rect 193364 142060 193370 142112
rect 146662 142032 146668 142044
rect 119816 142004 146668 142032
rect 114336 141992 114342 142004
rect 146662 141992 146668 142004
rect 146720 141992 146726 142044
rect 173250 141992 173256 142044
rect 173308 142032 173314 142044
rect 192110 142032 192116 142044
rect 173308 142004 192116 142032
rect 173308 141992 173314 142004
rect 192110 141992 192116 142004
rect 192168 141992 192174 142044
rect 119982 141924 119988 141976
rect 120040 141964 120046 141976
rect 151538 141964 151544 141976
rect 120040 141936 151544 141964
rect 120040 141924 120046 141936
rect 151538 141924 151544 141936
rect 151596 141924 151602 141976
rect 172422 141924 172428 141976
rect 172480 141964 172486 141976
rect 193398 141964 193404 141976
rect 172480 141936 193404 141964
rect 172480 141924 172486 141936
rect 193398 141924 193404 141936
rect 193456 141924 193462 141976
rect 105446 141856 105452 141908
rect 105504 141896 105510 141908
rect 138474 141896 138480 141908
rect 105504 141868 138480 141896
rect 105504 141856 105510 141868
rect 138474 141856 138480 141868
rect 138532 141856 138538 141908
rect 158346 141856 158352 141908
rect 158404 141896 158410 141908
rect 190730 141896 190736 141908
rect 158404 141868 190736 141896
rect 158404 141856 158410 141868
rect 190730 141856 190736 141868
rect 190788 141856 190794 141908
rect 115566 141788 115572 141840
rect 115624 141828 115630 141840
rect 148502 141828 148508 141840
rect 115624 141800 148508 141828
rect 115624 141788 115630 141800
rect 148502 141788 148508 141800
rect 148560 141788 148566 141840
rect 156506 141788 156512 141840
rect 156564 141828 156570 141840
rect 190638 141828 190644 141840
rect 156564 141800 190644 141828
rect 156564 141788 156570 141800
rect 190638 141788 190644 141800
rect 190696 141788 190702 141840
rect 118142 141720 118148 141772
rect 118200 141760 118206 141772
rect 152274 141760 152280 141772
rect 118200 141732 152280 141760
rect 118200 141720 118206 141732
rect 152274 141720 152280 141732
rect 152332 141720 152338 141772
rect 158622 141720 158628 141772
rect 158680 141760 158686 141772
rect 193766 141760 193772 141772
rect 158680 141732 193772 141760
rect 158680 141720 158686 141732
rect 193766 141720 193772 141732
rect 193824 141720 193830 141772
rect 115014 141652 115020 141704
rect 115072 141692 115078 141704
rect 149790 141692 149796 141704
rect 115072 141664 149796 141692
rect 115072 141652 115078 141664
rect 149790 141652 149796 141664
rect 149848 141652 149854 141704
rect 156966 141652 156972 141704
rect 157024 141692 157030 141704
rect 191190 141692 191196 141704
rect 157024 141664 191196 141692
rect 157024 141652 157030 141664
rect 191190 141652 191196 141664
rect 191248 141652 191254 141704
rect 113818 141584 113824 141636
rect 113876 141624 113882 141636
rect 148318 141624 148324 141636
rect 113876 141596 148324 141624
rect 113876 141584 113882 141596
rect 148318 141584 148324 141596
rect 148376 141584 148382 141636
rect 153102 141584 153108 141636
rect 153160 141624 153166 141636
rect 191098 141624 191104 141636
rect 153160 141596 191104 141624
rect 153160 141584 153166 141596
rect 191098 141584 191104 141596
rect 191156 141584 191162 141636
rect 95970 141516 95976 141568
rect 96028 141556 96034 141568
rect 139946 141556 139952 141568
rect 96028 141528 139952 141556
rect 96028 141516 96034 141528
rect 139946 141516 139952 141528
rect 140004 141516 140010 141568
rect 165154 141516 165160 141568
rect 165212 141556 165218 141568
rect 206278 141556 206284 141568
rect 165212 141528 206284 141556
rect 165212 141516 165218 141528
rect 206278 141516 206284 141528
rect 206336 141516 206342 141568
rect 117866 141448 117872 141500
rect 117924 141488 117930 141500
rect 178126 141488 178132 141500
rect 117924 141460 178132 141488
rect 117924 141448 117930 141460
rect 178126 141448 178132 141460
rect 178184 141448 178190 141500
rect 190638 141448 190644 141500
rect 190696 141488 190702 141500
rect 395338 141488 395344 141500
rect 190696 141460 395344 141488
rect 190696 141448 190702 141460
rect 395338 141448 395344 141460
rect 395396 141448 395402 141500
rect 106734 141380 106740 141432
rect 106792 141420 106798 141432
rect 172514 141420 172520 141432
rect 106792 141392 172520 141420
rect 106792 141380 106798 141392
rect 172514 141380 172520 141392
rect 172572 141380 172578 141432
rect 174814 141380 174820 141432
rect 174872 141420 174878 141432
rect 190822 141420 190828 141432
rect 174872 141392 190828 141420
rect 174872 141380 174878 141392
rect 190822 141380 190828 141392
rect 190880 141380 190886 141432
rect 193306 141380 193312 141432
rect 193364 141420 193370 141432
rect 518894 141420 518900 141432
rect 193364 141392 518900 141420
rect 193364 141380 193370 141392
rect 518894 141380 518900 141392
rect 518952 141380 518958 141432
rect 3510 141312 3516 141364
rect 3568 141352 3574 141364
rect 8938 141352 8944 141364
rect 3568 141324 8944 141352
rect 3568 141312 3574 141324
rect 8938 141312 8944 141324
rect 8996 141312 9002 141364
rect 115658 141312 115664 141364
rect 115716 141352 115722 141364
rect 145558 141352 145564 141364
rect 115716 141324 145564 141352
rect 115716 141312 115722 141324
rect 145558 141312 145564 141324
rect 145616 141312 145622 141364
rect 174538 141312 174544 141364
rect 174596 141352 174602 141364
rect 190638 141352 190644 141364
rect 174596 141324 190644 141352
rect 174596 141312 174602 141324
rect 190638 141312 190644 141324
rect 190696 141312 190702 141364
rect 119614 140836 119620 140888
rect 119672 140876 119678 140888
rect 119890 140876 119896 140888
rect 119672 140848 119896 140876
rect 119672 140836 119678 140848
rect 119890 140836 119896 140848
rect 119948 140836 119954 140888
rect 4798 140768 4804 140820
rect 4856 140808 4862 140820
rect 158346 140808 158352 140820
rect 4856 140780 158352 140808
rect 4856 140768 4862 140780
rect 158346 140768 158352 140780
rect 158404 140768 158410 140820
rect 147858 140740 147864 140752
rect 118666 140712 147864 140740
rect 117130 140632 117136 140684
rect 117188 140672 117194 140684
rect 118666 140672 118694 140712
rect 147858 140700 147864 140712
rect 147916 140700 147922 140752
rect 151906 140700 151912 140752
rect 151964 140740 151970 140752
rect 152550 140740 152556 140752
rect 151964 140712 152556 140740
rect 151964 140700 151970 140712
rect 152550 140700 152556 140712
rect 152608 140700 152614 140752
rect 164326 140700 164332 140752
rect 164384 140740 164390 140752
rect 164970 140740 164976 140752
rect 164384 140712 164976 140740
rect 164384 140700 164390 140712
rect 164970 140700 164976 140712
rect 165028 140700 165034 140752
rect 182818 140700 182824 140752
rect 182876 140740 182882 140752
rect 192386 140740 192392 140752
rect 182876 140712 192392 140740
rect 182876 140700 182882 140712
rect 192386 140700 192392 140712
rect 192444 140700 192450 140752
rect 117188 140644 118694 140672
rect 117188 140632 117194 140644
rect 119246 140632 119252 140684
rect 119304 140672 119310 140684
rect 123202 140672 123208 140684
rect 119304 140644 123208 140672
rect 119304 140632 119310 140644
rect 123202 140632 123208 140644
rect 123260 140632 123266 140684
rect 185946 140632 185952 140684
rect 186004 140672 186010 140684
rect 190730 140672 190736 140684
rect 186004 140644 190736 140672
rect 186004 140632 186010 140644
rect 190730 140632 190736 140644
rect 190788 140632 190794 140684
rect 114002 140564 114008 140616
rect 114060 140604 114066 140616
rect 124858 140604 124864 140616
rect 114060 140576 124864 140604
rect 114060 140564 114066 140576
rect 124858 140564 124864 140576
rect 124916 140564 124922 140616
rect 180150 140564 180156 140616
rect 180208 140604 180214 140616
rect 196710 140604 196716 140616
rect 180208 140576 196716 140604
rect 180208 140564 180214 140576
rect 196710 140564 196716 140576
rect 196768 140564 196774 140616
rect 115842 140496 115848 140548
rect 115900 140536 115906 140548
rect 132034 140536 132040 140548
rect 115900 140508 132040 140536
rect 115900 140496 115906 140508
rect 132034 140496 132040 140508
rect 132092 140496 132098 140548
rect 178678 140496 178684 140548
rect 178736 140536 178742 140548
rect 195330 140536 195336 140548
rect 178736 140508 195336 140536
rect 178736 140496 178742 140508
rect 195330 140496 195336 140508
rect 195388 140496 195394 140548
rect 112530 140428 112536 140480
rect 112588 140468 112594 140480
rect 131850 140468 131856 140480
rect 112588 140440 131856 140468
rect 112588 140428 112594 140440
rect 131850 140428 131856 140440
rect 131908 140428 131914 140480
rect 180058 140428 180064 140480
rect 180116 140468 180122 140480
rect 199102 140468 199108 140480
rect 180116 140440 199108 140468
rect 180116 140428 180122 140440
rect 199102 140428 199108 140440
rect 199160 140428 199166 140480
rect 110874 140360 110880 140412
rect 110932 140400 110938 140412
rect 131942 140400 131948 140412
rect 110932 140372 131948 140400
rect 110932 140360 110938 140372
rect 131942 140360 131948 140372
rect 132000 140360 132006 140412
rect 178770 140360 178776 140412
rect 178828 140400 178834 140412
rect 197814 140400 197820 140412
rect 178828 140372 197820 140400
rect 178828 140360 178834 140372
rect 197814 140360 197820 140372
rect 197872 140360 197878 140412
rect 102778 140292 102784 140344
rect 102836 140332 102842 140344
rect 133138 140332 133144 140344
rect 102836 140304 133144 140332
rect 102836 140292 102842 140304
rect 133138 140292 133144 140304
rect 133196 140292 133202 140344
rect 173158 140292 173164 140344
rect 173216 140332 173222 140344
rect 193490 140332 193496 140344
rect 173216 140304 193496 140332
rect 173216 140292 173222 140304
rect 193490 140292 193496 140304
rect 193548 140292 193554 140344
rect 113910 140224 113916 140276
rect 113968 140264 113974 140276
rect 145466 140264 145472 140276
rect 113968 140236 145472 140264
rect 113968 140224 113974 140236
rect 145466 140224 145472 140236
rect 145524 140224 145530 140276
rect 163774 140224 163780 140276
rect 163832 140264 163838 140276
rect 186314 140264 186320 140276
rect 163832 140236 186320 140264
rect 163832 140224 163838 140236
rect 186314 140224 186320 140236
rect 186372 140224 186378 140276
rect 123478 140156 123484 140208
rect 123536 140196 123542 140208
rect 149606 140196 149612 140208
rect 123536 140168 149612 140196
rect 123536 140156 123542 140168
rect 149606 140156 149612 140168
rect 149664 140156 149670 140208
rect 169938 140156 169944 140208
rect 169996 140196 170002 140208
rect 204898 140196 204904 140208
rect 169996 140168 204904 140196
rect 169996 140156 170002 140168
rect 204898 140156 204904 140168
rect 204956 140156 204962 140208
rect 103974 140088 103980 140140
rect 104032 140128 104038 140140
rect 137186 140128 137192 140140
rect 104032 140100 137192 140128
rect 104032 140088 104038 140100
rect 137186 140088 137192 140100
rect 137244 140088 137250 140140
rect 154666 140088 154672 140140
rect 154724 140128 154730 140140
rect 214742 140128 214748 140140
rect 154724 140100 214748 140128
rect 154724 140088 154730 140100
rect 214742 140088 214748 140100
rect 214800 140088 214806 140140
rect 97166 140020 97172 140072
rect 97224 140060 97230 140072
rect 138382 140060 138388 140072
rect 97224 140032 138388 140060
rect 97224 140020 97230 140032
rect 138382 140020 138388 140032
rect 138440 140020 138446 140072
rect 155770 140020 155776 140072
rect 155828 140060 155834 140072
rect 189534 140060 189540 140072
rect 155828 140032 189540 140060
rect 155828 140020 155834 140032
rect 189534 140020 189540 140032
rect 189592 140020 189598 140072
rect 193582 140020 193588 140072
rect 193640 140060 193646 140072
rect 335354 140060 335360 140072
rect 193640 140032 335360 140060
rect 193640 140020 193646 140032
rect 335354 140020 335360 140032
rect 335412 140020 335418 140072
rect 116670 139952 116676 140004
rect 116728 139992 116734 140004
rect 123478 139992 123484 140004
rect 116728 139964 123484 139992
rect 116728 139952 116734 139964
rect 123478 139952 123484 139964
rect 123536 139952 123542 140004
rect 146662 139952 146668 140004
rect 146720 139992 146726 140004
rect 146938 139992 146944 140004
rect 146720 139964 146944 139992
rect 146720 139952 146726 139964
rect 146938 139952 146944 139964
rect 146996 139952 147002 140004
rect 185578 139952 185584 140004
rect 185636 139992 185642 140004
rect 190454 139992 190460 140004
rect 185636 139964 190460 139992
rect 185636 139952 185642 139964
rect 190454 139952 190460 139964
rect 190512 139952 190518 140004
rect 185854 139884 185860 139936
rect 185912 139924 185918 139936
rect 193582 139924 193588 139936
rect 185912 139896 193588 139924
rect 185912 139884 185918 139896
rect 193582 139884 193588 139896
rect 193640 139884 193646 139936
rect 188338 139816 188344 139868
rect 188396 139856 188402 139868
rect 188890 139856 188896 139868
rect 188396 139828 188896 139856
rect 188396 139816 188402 139828
rect 188890 139816 188896 139828
rect 188948 139816 188954 139868
rect 119798 139544 119804 139596
rect 119856 139584 119862 139596
rect 124950 139584 124956 139596
rect 119856 139556 124956 139584
rect 119856 139544 119862 139556
rect 124950 139544 124956 139556
rect 125008 139544 125014 139596
rect 214742 139408 214748 139460
rect 214800 139448 214806 139460
rect 580442 139448 580448 139460
rect 214800 139420 580448 139448
rect 214800 139408 214806 139420
rect 580442 139408 580448 139420
rect 580500 139408 580506 139460
rect 128998 139312 129004 139324
rect 118666 139284 129004 139312
rect 116762 138660 116768 138712
rect 116820 138700 116826 138712
rect 118666 138700 118694 139284
rect 128998 139272 129004 139284
rect 129056 139272 129062 139324
rect 170582 139272 170588 139324
rect 170640 139272 170646 139324
rect 188246 139272 188252 139324
rect 188304 139272 188310 139324
rect 170600 138768 170628 139272
rect 188264 138836 188292 139272
rect 192754 138864 192760 138916
rect 192812 138904 192818 138916
rect 202230 138904 202236 138916
rect 192812 138876 202236 138904
rect 192812 138864 192818 138876
rect 202230 138864 202236 138876
rect 202288 138864 202294 138916
rect 205082 138836 205088 138848
rect 180766 138808 186314 138836
rect 188264 138808 205088 138836
rect 180766 138768 180794 138808
rect 170600 138740 180794 138768
rect 186286 138768 186314 138808
rect 205082 138796 205088 138808
rect 205140 138796 205146 138848
rect 196434 138768 196440 138780
rect 186286 138740 196440 138768
rect 196434 138728 196440 138740
rect 196492 138728 196498 138780
rect 116820 138672 118694 138700
rect 116820 138660 116826 138672
rect 188982 138660 188988 138712
rect 189040 138700 189046 138712
rect 580626 138700 580632 138712
rect 189040 138672 580632 138700
rect 189040 138660 189046 138672
rect 580626 138660 580632 138672
rect 580684 138660 580690 138712
rect 188982 137776 188988 137828
rect 189040 137816 189046 137828
rect 197538 137816 197544 137828
rect 189040 137788 197544 137816
rect 189040 137776 189046 137788
rect 197538 137776 197544 137788
rect 197596 137776 197602 137828
rect 200850 137096 200856 137148
rect 200908 137136 200914 137148
rect 203702 137136 203708 137148
rect 200908 137108 203708 137136
rect 200908 137096 200914 137108
rect 203702 137096 203708 137108
rect 203760 137096 203766 137148
rect 3418 136620 3424 136672
rect 3476 136660 3482 136672
rect 105354 136660 105360 136672
rect 3476 136632 105360 136660
rect 3476 136620 3482 136632
rect 105354 136620 105360 136632
rect 105412 136660 105418 136672
rect 108114 136660 108120 136672
rect 105412 136632 108120 136660
rect 105412 136620 105418 136632
rect 108114 136620 108120 136632
rect 108172 136620 108178 136672
rect 203702 136620 203708 136672
rect 203760 136660 203766 136672
rect 580166 136660 580172 136672
rect 203760 136632 580172 136660
rect 203760 136620 203766 136632
rect 580166 136620 580172 136632
rect 580224 136620 580230 136672
rect 118234 135872 118240 135924
rect 118292 135912 118298 135924
rect 119982 135912 119988 135924
rect 118292 135884 119988 135912
rect 118292 135872 118298 135884
rect 119982 135872 119988 135884
rect 120040 135872 120046 135924
rect 196618 124856 196624 124908
rect 196676 124896 196682 124908
rect 206462 124896 206468 124908
rect 196676 124868 206468 124896
rect 196676 124856 196682 124868
rect 206462 124856 206468 124868
rect 206520 124856 206526 124908
rect 206462 124176 206468 124228
rect 206520 124216 206526 124228
rect 580166 124216 580172 124228
rect 206520 124188 580172 124216
rect 206520 124176 206526 124188
rect 580166 124176 580172 124188
rect 580224 124176 580230 124228
rect 3142 121388 3148 121440
rect 3200 121428 3206 121440
rect 106734 121428 106740 121440
rect 3200 121400 106740 121428
rect 3200 121388 3206 121400
rect 106734 121388 106740 121400
rect 106792 121388 106798 121440
rect 3234 117240 3240 117292
rect 3292 117280 3298 117292
rect 103974 117280 103980 117292
rect 3292 117252 103980 117280
rect 3292 117240 3298 117252
rect 103974 117240 103980 117252
rect 104032 117240 104038 117292
rect 210602 112412 210608 112464
rect 210660 112452 210666 112464
rect 580166 112452 580172 112464
rect 210660 112424 580172 112452
rect 210660 112412 210666 112424
rect 580166 112412 580172 112424
rect 580224 112412 580230 112464
rect 3418 111800 3424 111852
rect 3476 111840 3482 111852
rect 113634 111840 113640 111852
rect 3476 111812 113640 111840
rect 3476 111800 3482 111812
rect 113634 111800 113640 111812
rect 113692 111800 113698 111852
rect 3418 108944 3424 108996
rect 3476 108984 3482 108996
rect 102134 108984 102140 108996
rect 3476 108956 102140 108984
rect 3476 108944 3482 108956
rect 102134 108944 102140 108956
rect 102192 108984 102198 108996
rect 102594 108984 102600 108996
rect 102192 108956 102600 108984
rect 102192 108944 102198 108956
rect 102594 108944 102600 108956
rect 102652 108944 102658 108996
rect 102134 108264 102140 108316
rect 102192 108304 102198 108316
rect 112254 108304 112260 108316
rect 102192 108276 112260 108304
rect 102192 108264 102198 108276
rect 112254 108264 112260 108276
rect 112312 108264 112318 108316
rect 194042 105408 194048 105460
rect 194100 105448 194106 105460
rect 202322 105448 202328 105460
rect 194100 105420 202328 105448
rect 194100 105408 194106 105420
rect 202322 105408 202328 105420
rect 202380 105408 202386 105460
rect 3418 103504 3424 103556
rect 3476 103544 3482 103556
rect 119154 103544 119160 103556
rect 3476 103516 119160 103544
rect 3476 103504 3482 103516
rect 119154 103504 119160 103516
rect 119212 103504 119218 103556
rect 3418 96636 3424 96688
rect 3476 96676 3482 96688
rect 117774 96676 117780 96688
rect 3476 96648 117780 96676
rect 3476 96636 3482 96648
rect 117774 96636 117780 96648
rect 117832 96636 117838 96688
rect 119338 95140 119344 95192
rect 119396 95180 119402 95192
rect 120534 95180 120540 95192
rect 119396 95152 120540 95180
rect 119396 95140 119402 95152
rect 120534 95140 120540 95152
rect 120592 95140 120598 95192
rect 3142 93780 3148 93832
rect 3200 93820 3206 93832
rect 115014 93820 115020 93832
rect 3200 93792 115020 93820
rect 3200 93780 3206 93792
rect 115014 93780 115020 93792
rect 115072 93780 115078 93832
rect 115014 92488 115020 92540
rect 115072 92528 115078 92540
rect 119338 92528 119344 92540
rect 115072 92500 119344 92528
rect 115072 92488 115078 92500
rect 119338 92488 119344 92500
rect 119396 92488 119402 92540
rect 191282 91060 191288 91112
rect 191340 91100 191346 91112
rect 198182 91100 198188 91112
rect 191340 91072 198188 91100
rect 191340 91060 191346 91072
rect 198182 91060 198188 91072
rect 198240 91060 198246 91112
rect 189718 85144 189724 85196
rect 189776 85144 189782 85196
rect 189736 84924 189764 85144
rect 189718 84872 189724 84924
rect 189776 84872 189782 84924
rect 189166 84804 189172 84856
rect 189224 84844 189230 84856
rect 189626 84844 189632 84856
rect 189224 84816 189632 84844
rect 189224 84804 189230 84816
rect 189626 84804 189632 84816
rect 189684 84804 189690 84856
rect 3418 84192 3424 84244
rect 3476 84232 3482 84244
rect 98546 84232 98552 84244
rect 3476 84204 98552 84232
rect 3476 84192 3482 84204
rect 98546 84192 98552 84204
rect 98604 84192 98610 84244
rect 189166 82084 189172 82136
rect 189224 82124 189230 82136
rect 206462 82124 206468 82136
rect 189224 82096 206468 82124
rect 189224 82084 189230 82096
rect 206462 82084 206468 82096
rect 206520 82084 206526 82136
rect 188614 81676 188620 81728
rect 188672 81716 188678 81728
rect 188890 81716 188896 81728
rect 188672 81688 188896 81716
rect 188672 81676 188678 81688
rect 188890 81676 188896 81688
rect 188948 81676 188954 81728
rect 3418 81336 3424 81388
rect 3476 81376 3482 81388
rect 108298 81376 108304 81388
rect 3476 81348 108304 81376
rect 3476 81336 3482 81348
rect 108298 81336 108304 81348
rect 108356 81336 108362 81388
rect 194226 81104 194232 81116
rect 176626 81076 194232 81104
rect 176626 81036 176654 81076
rect 194226 81064 194232 81076
rect 194284 81064 194290 81116
rect 168346 81008 176654 81036
rect 133846 80940 138014 80968
rect 108298 80860 108304 80912
rect 108356 80900 108362 80912
rect 120074 80900 120080 80912
rect 108356 80872 120080 80900
rect 108356 80860 108362 80872
rect 120074 80860 120080 80872
rect 120132 80860 120138 80912
rect 120902 80860 120908 80912
rect 120960 80900 120966 80912
rect 133846 80900 133874 80940
rect 120960 80872 131896 80900
rect 120960 80860 120966 80872
rect 105630 80792 105636 80844
rect 105688 80832 105694 80844
rect 105688 80804 131804 80832
rect 105688 80792 105694 80804
rect 113542 80724 113548 80776
rect 113600 80764 113606 80776
rect 113600 80736 124214 80764
rect 113600 80724 113606 80736
rect 112346 80656 112352 80708
rect 112404 80696 112410 80708
rect 112404 80668 123524 80696
rect 112404 80656 112410 80668
rect 117958 80588 117964 80640
rect 118016 80628 118022 80640
rect 118016 80600 118694 80628
rect 118016 80588 118022 80600
rect 118666 80492 118694 80600
rect 123496 80560 123524 80668
rect 124186 80628 124214 80736
rect 131776 80708 131804 80804
rect 131868 80708 131896 80872
rect 132052 80872 133874 80900
rect 132052 80764 132080 80872
rect 135226 80804 136634 80832
rect 135226 80764 135254 80804
rect 131960 80736 132080 80764
rect 133846 80736 135254 80764
rect 131758 80656 131764 80708
rect 131816 80656 131822 80708
rect 131850 80656 131856 80708
rect 131908 80656 131914 80708
rect 131960 80628 131988 80736
rect 132034 80656 132040 80708
rect 132092 80696 132098 80708
rect 133846 80696 133874 80736
rect 132092 80668 133874 80696
rect 136606 80696 136634 80804
rect 137986 80764 138014 80940
rect 137986 80736 140774 80764
rect 140746 80696 140774 80736
rect 136606 80668 139164 80696
rect 140746 80668 147306 80696
rect 132092 80656 132098 80668
rect 124186 80600 131988 80628
rect 132788 80600 136634 80628
rect 132788 80560 132816 80600
rect 123496 80532 132816 80560
rect 133156 80532 134104 80560
rect 123570 80492 123576 80504
rect 118666 80464 123576 80492
rect 123570 80452 123576 80464
rect 123628 80452 123634 80504
rect 131758 80452 131764 80504
rect 131816 80492 131822 80504
rect 133156 80492 133184 80532
rect 131816 80464 133184 80492
rect 133340 80464 134012 80492
rect 131816 80452 131822 80464
rect 119614 80384 119620 80436
rect 119672 80424 119678 80436
rect 126238 80424 126244 80436
rect 119672 80396 126244 80424
rect 119672 80384 119678 80396
rect 126238 80384 126244 80396
rect 126296 80384 126302 80436
rect 119246 80316 119252 80368
rect 119304 80356 119310 80368
rect 126330 80356 126336 80368
rect 119304 80328 126336 80356
rect 119304 80316 119310 80328
rect 126330 80316 126336 80328
rect 126388 80316 126394 80368
rect 128446 80316 128452 80368
rect 128504 80356 128510 80368
rect 131850 80356 131856 80368
rect 128504 80328 131856 80356
rect 128504 80316 128510 80328
rect 131850 80316 131856 80328
rect 131908 80316 131914 80368
rect 133340 80356 133368 80464
rect 131960 80328 133368 80356
rect 133984 80356 134012 80464
rect 134076 80424 134104 80532
rect 136606 80492 136634 80600
rect 139136 80560 139164 80668
rect 139136 80532 140130 80560
rect 136606 80464 140038 80492
rect 134076 80396 139946 80424
rect 133984 80328 134610 80356
rect 128630 80248 128636 80300
rect 128688 80288 128694 80300
rect 131960 80288 131988 80328
rect 128688 80260 131988 80288
rect 128688 80248 128694 80260
rect 128538 80180 128544 80232
rect 128596 80220 128602 80232
rect 132218 80220 132224 80232
rect 128596 80192 132224 80220
rect 128596 80180 128602 80192
rect 132218 80180 132224 80192
rect 132276 80180 132282 80232
rect 134582 80220 134610 80328
rect 132328 80192 133368 80220
rect 134582 80192 138382 80220
rect 132034 80112 132040 80164
rect 132092 80152 132098 80164
rect 132328 80152 132356 80192
rect 132092 80124 132356 80152
rect 133340 80152 133368 80192
rect 133340 80124 134518 80152
rect 132092 80112 132098 80124
rect 126946 80056 132908 80084
rect 124582 79976 124588 80028
rect 124640 80016 124646 80028
rect 126946 80016 126974 80056
rect 132880 80016 132908 80056
rect 124640 79988 126974 80016
rect 129568 79988 132678 80016
rect 132880 79988 133046 80016
rect 124640 79976 124646 79988
rect 125226 79840 125232 79892
rect 125284 79880 125290 79892
rect 129568 79880 129596 79988
rect 132540 79908 132546 79960
rect 132598 79908 132604 79960
rect 132650 79948 132678 79988
rect 133018 79960 133046 79988
rect 133294 79988 134150 80016
rect 132908 79948 132914 79960
rect 132650 79920 132914 79948
rect 132908 79908 132914 79920
rect 132966 79908 132972 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 125284 79852 129596 79880
rect 125284 79840 125290 79852
rect 132558 79756 132586 79908
rect 133294 79880 133322 79988
rect 134122 79960 134150 79988
rect 134490 79960 134518 80124
rect 134582 79988 135806 80016
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133920 79908 133926 79960
rect 133978 79948 133984 79960
rect 134104 79948 134110 79960
rect 133978 79908 134012 79948
rect 132696 79852 133322 79880
rect 101214 79704 101220 79756
rect 101272 79744 101278 79756
rect 101272 79716 132494 79744
rect 132558 79716 132592 79756
rect 101272 79704 101278 79716
rect 97534 79636 97540 79688
rect 97592 79676 97598 79688
rect 128998 79676 129004 79688
rect 97592 79648 129004 79676
rect 97592 79636 97598 79648
rect 128998 79636 129004 79648
rect 129056 79636 129062 79688
rect 132466 79676 132494 79716
rect 132586 79704 132592 79716
rect 132644 79704 132650 79756
rect 132696 79676 132724 79852
rect 133276 79772 133282 79824
rect 133334 79772 133340 79824
rect 133294 79744 133322 79772
rect 132466 79648 132724 79676
rect 132880 79716 133322 79744
rect 115106 79568 115112 79620
rect 115164 79608 115170 79620
rect 122834 79608 122840 79620
rect 115164 79580 122840 79608
rect 115164 79568 115170 79580
rect 122834 79568 122840 79580
rect 122892 79568 122898 79620
rect 131298 79568 131304 79620
rect 131356 79608 131362 79620
rect 132880 79608 132908 79716
rect 133138 79636 133144 79688
rect 133196 79676 133202 79688
rect 133386 79676 133414 79908
rect 133828 79840 133834 79892
rect 133886 79840 133892 79892
rect 133552 79772 133558 79824
rect 133610 79772 133616 79824
rect 133644 79772 133650 79824
rect 133702 79772 133708 79824
rect 133570 79688 133598 79772
rect 133196 79648 133414 79676
rect 133196 79636 133202 79648
rect 133506 79636 133512 79688
rect 133564 79648 133598 79688
rect 133662 79688 133690 79772
rect 133662 79648 133696 79688
rect 133564 79636 133570 79648
rect 133690 79636 133696 79648
rect 133748 79636 133754 79688
rect 131356 79580 132908 79608
rect 133846 79608 133874 79840
rect 133984 79824 134012 79908
rect 134076 79908 134110 79948
rect 134162 79908 134168 79960
rect 134472 79908 134478 79960
rect 134530 79908 134536 79960
rect 133966 79772 133972 79824
rect 134024 79772 134030 79824
rect 133846 79580 133966 79608
rect 131356 79568 131362 79580
rect 113818 79500 113824 79552
rect 113876 79540 113882 79552
rect 127526 79540 127532 79552
rect 113876 79512 127532 79540
rect 113876 79500 113882 79512
rect 127526 79500 127532 79512
rect 127584 79500 127590 79552
rect 96062 79432 96068 79484
rect 96120 79472 96126 79484
rect 129274 79472 129280 79484
rect 96120 79444 129280 79472
rect 96120 79432 96126 79444
rect 129274 79432 129280 79444
rect 129332 79432 129338 79484
rect 121178 79364 121184 79416
rect 121236 79404 121242 79416
rect 133322 79404 133328 79416
rect 121236 79376 133328 79404
rect 121236 79364 121242 79376
rect 133322 79364 133328 79376
rect 133380 79364 133386 79416
rect 133782 79364 133788 79416
rect 133840 79404 133846 79416
rect 133938 79404 133966 79580
rect 133840 79376 133966 79404
rect 134076 79404 134104 79908
rect 134288 79840 134294 79892
rect 134346 79880 134352 79892
rect 134582 79880 134610 79988
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135484 79908 135490 79960
rect 135542 79908 135548 79960
rect 135668 79948 135674 79960
rect 135640 79908 135674 79948
rect 135726 79908 135732 79960
rect 134346 79852 134610 79880
rect 134346 79840 134352 79852
rect 134196 79772 134202 79824
rect 134254 79772 134260 79824
rect 134656 79812 134662 79824
rect 134444 79784 134662 79812
rect 134214 79688 134242 79772
rect 134444 79688 134472 79784
rect 134656 79772 134662 79784
rect 134714 79772 134720 79824
rect 134840 79772 134846 79824
rect 134898 79772 134904 79824
rect 135024 79812 135030 79824
rect 134996 79772 135030 79812
rect 135082 79772 135088 79824
rect 135208 79772 135214 79824
rect 135266 79772 135272 79824
rect 134150 79636 134156 79688
rect 134208 79648 134242 79688
rect 134208 79636 134214 79648
rect 134426 79636 134432 79688
rect 134484 79636 134490 79688
rect 134858 79608 134886 79772
rect 134996 79620 135024 79772
rect 135226 79688 135254 79772
rect 135410 79688 135438 79908
rect 135226 79648 135260 79688
rect 135254 79636 135260 79648
rect 135312 79636 135318 79688
rect 135346 79636 135352 79688
rect 135404 79648 135438 79688
rect 135404 79636 135410 79648
rect 134398 79580 134886 79608
rect 134242 79432 134248 79484
rect 134300 79472 134306 79484
rect 134398 79472 134426 79580
rect 134978 79568 134984 79620
rect 135036 79568 135042 79620
rect 134702 79500 134708 79552
rect 134760 79540 134766 79552
rect 135502 79540 135530 79908
rect 135640 79688 135668 79908
rect 135778 79880 135806 79988
rect 136882 79988 137278 80016
rect 136882 79960 136910 79988
rect 135944 79908 135950 79960
rect 136002 79948 136008 79960
rect 136002 79908 136036 79948
rect 136128 79908 136134 79960
rect 136186 79908 136192 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 136312 79908 136318 79960
rect 136370 79948 136376 79960
rect 136496 79948 136502 79960
rect 136370 79908 136404 79948
rect 135778 79852 135944 79880
rect 135916 79824 135944 79852
rect 135898 79772 135904 79824
rect 135956 79772 135962 79824
rect 136008 79688 136036 79908
rect 136146 79756 136174 79908
rect 136238 79880 136266 79908
rect 136238 79852 136312 79880
rect 136146 79716 136180 79756
rect 136174 79704 136180 79716
rect 136232 79704 136238 79756
rect 135622 79636 135628 79688
rect 135680 79636 135686 79688
rect 135990 79636 135996 79688
rect 136048 79636 136054 79688
rect 135898 79568 135904 79620
rect 135956 79608 135962 79620
rect 136284 79608 136312 79852
rect 136376 79620 136404 79908
rect 136468 79908 136502 79948
rect 136554 79908 136560 79960
rect 136864 79908 136870 79960
rect 136922 79908 136928 79960
rect 137048 79948 137054 79960
rect 137020 79908 137054 79948
rect 137106 79908 137112 79960
rect 136468 79688 136496 79908
rect 136450 79636 136456 79688
rect 136508 79636 136514 79688
rect 137020 79676 137048 79908
rect 137140 79880 137146 79892
rect 137112 79840 137146 79880
rect 137198 79840 137204 79892
rect 137112 79756 137140 79840
rect 137094 79704 137100 79756
rect 137152 79704 137158 79756
rect 136928 79648 137048 79676
rect 136928 79620 136956 79648
rect 135956 79580 136312 79608
rect 135956 79568 135962 79580
rect 136358 79568 136364 79620
rect 136416 79568 136422 79620
rect 136910 79568 136916 79620
rect 136968 79568 136974 79620
rect 137002 79568 137008 79620
rect 137060 79608 137066 79620
rect 137250 79608 137278 79988
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137784 79908 137790 79960
rect 137842 79908 137848 79960
rect 137876 79908 137882 79960
rect 137934 79908 137940 79960
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 137060 79580 137278 79608
rect 137060 79568 137066 79580
rect 137462 79568 137468 79620
rect 137520 79608 137526 79620
rect 137618 79608 137646 79908
rect 137520 79580 137646 79608
rect 137802 79620 137830 79908
rect 137894 79744 137922 79908
rect 138078 79880 138106 79908
rect 138032 79852 138106 79880
rect 137894 79716 137968 79744
rect 137940 79620 137968 79716
rect 138032 79620 138060 79852
rect 138170 79824 138198 79908
rect 138354 79892 138382 80192
rect 138538 79988 139348 80016
rect 138538 79892 138566 79988
rect 138704 79948 138710 79960
rect 138630 79920 138710 79948
rect 138336 79840 138342 79892
rect 138394 79840 138400 79892
rect 138520 79840 138526 79892
rect 138578 79840 138584 79892
rect 138106 79772 138112 79824
rect 138164 79784 138198 79824
rect 138164 79772 138170 79784
rect 138630 79688 138658 79920
rect 138704 79908 138710 79920
rect 138762 79908 138768 79960
rect 138980 79908 138986 79960
rect 139038 79948 139044 79960
rect 139038 79920 139210 79948
rect 139038 79908 139044 79920
rect 138796 79880 138802 79892
rect 138768 79840 138802 79880
rect 138854 79840 138860 79892
rect 138888 79840 138894 79892
rect 138946 79880 138952 79892
rect 138946 79840 138980 79880
rect 138768 79756 138796 79840
rect 138952 79756 138980 79840
rect 139072 79772 139078 79824
rect 139130 79772 139136 79824
rect 138750 79704 138756 79756
rect 138808 79704 138814 79756
rect 138934 79704 138940 79756
rect 138992 79704 138998 79756
rect 139090 79688 139118 79772
rect 138566 79636 138572 79688
rect 138624 79648 138658 79688
rect 138624 79636 138630 79648
rect 139026 79636 139032 79688
rect 139084 79648 139118 79688
rect 139084 79636 139090 79648
rect 137802 79580 137836 79620
rect 137520 79568 137526 79580
rect 137830 79568 137836 79580
rect 137888 79568 137894 79620
rect 137922 79568 137928 79620
rect 137980 79568 137986 79620
rect 138014 79568 138020 79620
rect 138072 79568 138078 79620
rect 138842 79568 138848 79620
rect 138900 79608 138906 79620
rect 139182 79608 139210 79920
rect 138900 79580 139210 79608
rect 139320 79608 139348 79988
rect 139918 79960 139946 80396
rect 140010 80016 140038 80464
rect 140102 80356 140130 80532
rect 140102 80328 140222 80356
rect 140194 80084 140222 80328
rect 140194 80056 141648 80084
rect 140010 79988 141418 80016
rect 139532 79948 139538 79960
rect 139412 79920 139538 79948
rect 139412 79688 139440 79920
rect 139532 79908 139538 79920
rect 139590 79908 139596 79960
rect 139900 79908 139906 79960
rect 139958 79908 139964 79960
rect 139992 79908 139998 79960
rect 140050 79908 140056 79960
rect 141096 79948 141102 79960
rect 141068 79908 141102 79948
rect 141154 79908 141160 79960
rect 140010 79880 140038 79908
rect 139504 79852 140038 79880
rect 139504 79756 139532 79852
rect 140544 79840 140550 79892
rect 140602 79840 140608 79892
rect 140820 79840 140826 79892
rect 140878 79840 140884 79892
rect 140038 79772 140044 79824
rect 140096 79812 140102 79824
rect 140562 79812 140590 79840
rect 140096 79784 140590 79812
rect 140096 79772 140102 79784
rect 139486 79704 139492 79756
rect 139544 79704 139550 79756
rect 140838 79688 140866 79840
rect 141068 79688 141096 79908
rect 141188 79880 141194 79892
rect 141160 79840 141194 79880
rect 141246 79840 141252 79892
rect 141280 79840 141286 79892
rect 141338 79840 141344 79892
rect 141390 79880 141418 79988
rect 141620 79960 141648 80056
rect 141758 79988 144730 80016
rect 141620 79920 141654 79960
rect 141648 79908 141654 79920
rect 141706 79908 141712 79960
rect 141758 79880 141786 79988
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142108 79908 142114 79960
rect 142166 79908 142172 79960
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 142476 79908 142482 79960
rect 142534 79948 142540 79960
rect 142534 79920 142890 79948
rect 142534 79908 142540 79920
rect 141390 79852 141786 79880
rect 141832 79840 141838 79892
rect 141890 79840 141896 79892
rect 141160 79756 141188 79840
rect 141142 79704 141148 79756
rect 141200 79704 141206 79756
rect 141298 79688 141326 79840
rect 141464 79812 141470 79824
rect 141436 79772 141470 79812
rect 141522 79772 141528 79824
rect 141556 79772 141562 79824
rect 141614 79772 141620 79824
rect 141850 79812 141878 79840
rect 141712 79784 141878 79812
rect 141436 79688 141464 79772
rect 141574 79744 141602 79772
rect 141528 79716 141602 79744
rect 141528 79688 141556 79716
rect 139394 79636 139400 79688
rect 139452 79636 139458 79688
rect 140774 79636 140780 79688
rect 140832 79648 140866 79688
rect 140832 79636 140838 79648
rect 141050 79636 141056 79688
rect 141108 79636 141114 79688
rect 141298 79648 141332 79688
rect 141326 79636 141332 79648
rect 141384 79636 141390 79688
rect 141418 79636 141424 79688
rect 141476 79636 141482 79688
rect 141510 79636 141516 79688
rect 141568 79636 141574 79688
rect 141602 79636 141608 79688
rect 141660 79676 141666 79688
rect 141712 79676 141740 79784
rect 141942 79756 141970 79908
rect 141878 79704 141884 79756
rect 141936 79716 141970 79756
rect 141936 79704 141942 79716
rect 141660 79648 141740 79676
rect 141660 79636 141666 79648
rect 140406 79608 140412 79620
rect 139320 79580 140412 79608
rect 138900 79568 138906 79580
rect 140406 79568 140412 79580
rect 140464 79568 140470 79620
rect 142126 79608 142154 79908
rect 142402 79744 142430 79908
rect 142752 79840 142758 79892
rect 142810 79840 142816 79892
rect 142568 79812 142574 79824
rect 142540 79772 142574 79812
rect 142626 79772 142632 79824
rect 142402 79716 142476 79744
rect 142448 79688 142476 79716
rect 142540 79688 142568 79772
rect 142770 79744 142798 79840
rect 142632 79716 142798 79744
rect 142632 79688 142660 79716
rect 142430 79636 142436 79688
rect 142488 79636 142494 79688
rect 142522 79636 142528 79688
rect 142580 79636 142586 79688
rect 142614 79636 142620 79688
rect 142672 79636 142678 79688
rect 142246 79608 142252 79620
rect 142126 79580 142252 79608
rect 142246 79568 142252 79580
rect 142304 79568 142310 79620
rect 142862 79608 142890 79920
rect 143120 79908 143126 79960
rect 143178 79908 143184 79960
rect 143396 79908 143402 79960
rect 143454 79908 143460 79960
rect 144132 79948 144138 79960
rect 143552 79920 144138 79948
rect 143138 79688 143166 79908
rect 143074 79636 143080 79688
rect 143132 79648 143166 79688
rect 143132 79636 143138 79648
rect 143414 79620 143442 79908
rect 142816 79580 142890 79608
rect 142816 79552 142844 79580
rect 143350 79568 143356 79620
rect 143408 79580 143442 79620
rect 143408 79568 143414 79580
rect 143552 79552 143580 79920
rect 144132 79908 144138 79920
rect 144190 79908 144196 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 143672 79880 143678 79892
rect 143644 79840 143678 79880
rect 143730 79840 143736 79892
rect 143764 79840 143770 79892
rect 143822 79840 143828 79892
rect 143948 79840 143954 79892
rect 144006 79840 144012 79892
rect 144040 79840 144046 79892
rect 144098 79840 144104 79892
rect 143644 79688 143672 79840
rect 143626 79636 143632 79688
rect 143684 79636 143690 79688
rect 143782 79552 143810 79840
rect 143966 79620 143994 79840
rect 143902 79568 143908 79620
rect 143960 79580 143994 79620
rect 143960 79568 143966 79580
rect 144058 79552 144086 79840
rect 144242 79756 144270 79908
rect 144178 79704 144184 79756
rect 144236 79716 144270 79756
rect 144236 79704 144242 79716
rect 144178 79568 144184 79620
rect 144236 79608 144242 79620
rect 144334 79608 144362 79908
rect 144500 79840 144506 79892
rect 144558 79840 144564 79892
rect 144592 79840 144598 79892
rect 144650 79840 144656 79892
rect 144518 79688 144546 79840
rect 144454 79636 144460 79688
rect 144512 79648 144546 79688
rect 144512 79636 144518 79648
rect 144610 79620 144638 79840
rect 144236 79580 144362 79608
rect 144236 79568 144242 79580
rect 144546 79568 144552 79620
rect 144604 79580 144638 79620
rect 144702 79608 144730 79988
rect 147278 79960 147306 80668
rect 168346 80628 168374 81008
rect 188614 80996 188620 81048
rect 188672 81036 188678 81048
rect 202874 81036 202880 81048
rect 188672 81008 202880 81036
rect 188672 80996 188678 81008
rect 202874 80996 202880 81008
rect 202932 80996 202938 81048
rect 203702 80968 203708 80980
rect 177868 80940 203708 80968
rect 177868 80708 177896 80940
rect 203702 80928 203708 80940
rect 203760 80928 203766 80980
rect 207382 80900 207388 80912
rect 178006 80872 207388 80900
rect 178006 80708 178034 80872
rect 207382 80860 207388 80872
rect 207440 80860 207446 80912
rect 195330 80764 195336 80776
rect 177850 80656 177856 80708
rect 177908 80656 177914 80708
rect 177942 80656 177948 80708
rect 178000 80668 178034 80708
rect 178420 80736 195336 80764
rect 178000 80656 178006 80668
rect 178420 80628 178448 80736
rect 195330 80724 195336 80736
rect 195388 80724 195394 80776
rect 182818 80656 182824 80708
rect 182876 80696 182882 80708
rect 211982 80696 211988 80708
rect 182876 80668 211988 80696
rect 182876 80656 182882 80668
rect 211982 80656 211988 80668
rect 212040 80656 212046 80708
rect 159882 80600 168374 80628
rect 169634 80600 178448 80628
rect 151832 80056 152918 80084
rect 147462 79988 149882 80016
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 144960 79908 144966 79960
rect 145018 79908 145024 79960
rect 145052 79908 145058 79960
rect 145110 79908 145116 79960
rect 145144 79908 145150 79960
rect 145202 79908 145208 79960
rect 145420 79908 145426 79960
rect 145478 79908 145484 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 145972 79908 145978 79960
rect 146030 79908 146036 79960
rect 146064 79908 146070 79960
rect 146122 79908 146128 79960
rect 146432 79948 146438 79960
rect 146404 79908 146438 79948
rect 146490 79908 146496 79960
rect 146616 79908 146622 79960
rect 146674 79908 146680 79960
rect 146892 79908 146898 79960
rect 146950 79908 146956 79960
rect 147260 79908 147266 79960
rect 147318 79908 147324 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 144886 79824 144914 79908
rect 144822 79772 144828 79824
rect 144880 79784 144914 79824
rect 144880 79772 144886 79784
rect 144978 79756 145006 79908
rect 145070 79824 145098 79908
rect 145162 79880 145190 79908
rect 145162 79852 145236 79880
rect 145208 79824 145236 79852
rect 145070 79784 145104 79824
rect 145098 79772 145104 79784
rect 145156 79772 145162 79824
rect 145190 79772 145196 79824
rect 145248 79772 145254 79824
rect 144914 79704 144920 79756
rect 144972 79716 145006 79756
rect 144972 79704 144978 79716
rect 145006 79636 145012 79688
rect 145064 79676 145070 79688
rect 145438 79676 145466 79908
rect 145696 79880 145702 79892
rect 145668 79840 145702 79880
rect 145754 79840 145760 79892
rect 145668 79756 145696 79840
rect 145806 79756 145834 79908
rect 145990 79756 146018 79908
rect 145650 79704 145656 79756
rect 145708 79704 145714 79756
rect 145742 79704 145748 79756
rect 145800 79716 145834 79756
rect 145800 79704 145806 79716
rect 145926 79704 145932 79756
rect 145984 79716 146018 79756
rect 146082 79756 146110 79908
rect 146248 79880 146254 79892
rect 146220 79840 146254 79880
rect 146306 79840 146312 79892
rect 146220 79756 146248 79840
rect 146404 79756 146432 79908
rect 146082 79716 146116 79756
rect 145984 79704 145990 79716
rect 146110 79704 146116 79716
rect 146168 79704 146174 79756
rect 146202 79704 146208 79756
rect 146260 79704 146266 79756
rect 146386 79704 146392 79756
rect 146444 79704 146450 79756
rect 145064 79648 145466 79676
rect 145064 79636 145070 79648
rect 146018 79636 146024 79688
rect 146076 79676 146082 79688
rect 146634 79676 146662 79908
rect 146800 79840 146806 79892
rect 146858 79840 146864 79892
rect 146076 79648 146662 79676
rect 146076 79636 146082 79648
rect 145558 79608 145564 79620
rect 144702 79580 145564 79608
rect 144604 79568 144610 79580
rect 145558 79568 145564 79580
rect 145616 79568 145622 79620
rect 134760 79512 135530 79540
rect 134760 79500 134766 79512
rect 136726 79500 136732 79552
rect 136784 79540 136790 79552
rect 136784 79512 141096 79540
rect 136784 79500 136790 79512
rect 134300 79444 134426 79472
rect 134300 79432 134306 79444
rect 134886 79432 134892 79484
rect 134944 79472 134950 79484
rect 140774 79472 140780 79484
rect 134944 79444 140780 79472
rect 134944 79432 134950 79444
rect 140774 79432 140780 79444
rect 140832 79432 140838 79484
rect 141068 79472 141096 79512
rect 142798 79500 142804 79552
rect 142856 79500 142862 79552
rect 143534 79500 143540 79552
rect 143592 79500 143598 79552
rect 143782 79512 143816 79552
rect 143810 79500 143816 79512
rect 143868 79500 143874 79552
rect 144058 79512 144092 79552
rect 144086 79500 144092 79512
rect 144144 79500 144150 79552
rect 145466 79500 145472 79552
rect 145524 79540 145530 79552
rect 145834 79540 145840 79552
rect 145524 79512 145840 79540
rect 145524 79500 145530 79512
rect 145834 79500 145840 79512
rect 145892 79500 145898 79552
rect 146662 79500 146668 79552
rect 146720 79540 146726 79552
rect 146818 79540 146846 79840
rect 146910 79688 146938 79908
rect 147370 79824 147398 79908
rect 147306 79772 147312 79824
rect 147364 79784 147398 79824
rect 147364 79772 147370 79784
rect 147462 79756 147490 79988
rect 149854 79960 149882 79988
rect 150590 79988 151354 80016
rect 147536 79908 147542 79960
rect 147594 79908 147600 79960
rect 147720 79948 147726 79960
rect 147692 79908 147726 79948
rect 147778 79908 147784 79960
rect 148456 79908 148462 79960
rect 148514 79908 148520 79960
rect 148732 79908 148738 79960
rect 148790 79908 148796 79960
rect 148916 79908 148922 79960
rect 148974 79948 148980 79960
rect 148974 79908 149008 79948
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 149376 79908 149382 79960
rect 149434 79948 149440 79960
rect 149434 79908 149468 79948
rect 149652 79908 149658 79960
rect 149710 79908 149716 79960
rect 149836 79908 149842 79960
rect 149894 79908 149900 79960
rect 149928 79908 149934 79960
rect 149986 79908 149992 79960
rect 150480 79908 150486 79960
rect 150538 79908 150544 79960
rect 147398 79704 147404 79756
rect 147456 79716 147490 79756
rect 147456 79704 147462 79716
rect 147554 79688 147582 79908
rect 147692 79824 147720 79908
rect 147904 79840 147910 79892
rect 147962 79840 147968 79892
rect 148088 79840 148094 79892
rect 148146 79840 148152 79892
rect 148180 79840 148186 79892
rect 148238 79840 148244 79892
rect 147674 79772 147680 79824
rect 147732 79772 147738 79824
rect 146910 79648 146944 79688
rect 146938 79636 146944 79648
rect 146996 79636 147002 79688
rect 147490 79636 147496 79688
rect 147548 79648 147582 79688
rect 147548 79636 147554 79648
rect 147922 79620 147950 79840
rect 147922 79580 147956 79620
rect 147950 79568 147956 79580
rect 148008 79568 148014 79620
rect 146720 79512 146846 79540
rect 148106 79540 148134 79840
rect 148198 79688 148226 79840
rect 148364 79772 148370 79824
rect 148422 79772 148428 79824
rect 148198 79648 148232 79688
rect 148226 79636 148232 79648
rect 148284 79636 148290 79688
rect 148382 79608 148410 79772
rect 148474 79688 148502 79908
rect 148474 79648 148508 79688
rect 148502 79636 148508 79648
rect 148560 79636 148566 79688
rect 148594 79636 148600 79688
rect 148652 79676 148658 79688
rect 148750 79676 148778 79908
rect 148824 79840 148830 79892
rect 148882 79880 148888 79892
rect 148882 79840 148916 79880
rect 148888 79688 148916 79840
rect 148652 79648 148778 79676
rect 148652 79636 148658 79648
rect 148870 79636 148876 79688
rect 148928 79636 148934 79688
rect 148980 79608 149008 79908
rect 149210 79676 149238 79908
rect 149440 79688 149468 79908
rect 149560 79880 149566 79892
rect 149532 79840 149566 79880
rect 149618 79840 149624 79892
rect 149164 79648 149238 79676
rect 149054 79608 149060 79620
rect 148382 79580 148916 79608
rect 148980 79580 149060 79608
rect 148226 79540 148232 79552
rect 148106 79512 148232 79540
rect 146720 79500 146726 79512
rect 148226 79500 148232 79512
rect 148284 79500 148290 79552
rect 148888 79540 148916 79580
rect 149054 79568 149060 79580
rect 149112 79568 149118 79620
rect 148962 79540 148968 79552
rect 148888 79512 148968 79540
rect 148962 79500 148968 79512
rect 149020 79500 149026 79552
rect 149164 79540 149192 79648
rect 149422 79636 149428 79688
rect 149480 79636 149486 79688
rect 149238 79568 149244 79620
rect 149296 79608 149302 79620
rect 149532 79608 149560 79840
rect 149670 79688 149698 79908
rect 149606 79636 149612 79688
rect 149664 79648 149698 79688
rect 149664 79636 149670 79648
rect 149296 79580 149560 79608
rect 149296 79568 149302 79580
rect 149790 79568 149796 79620
rect 149848 79608 149854 79620
rect 149946 79608 149974 79908
rect 150296 79840 150302 79892
rect 150354 79840 150360 79892
rect 150314 79756 150342 79840
rect 150498 79756 150526 79908
rect 150250 79704 150256 79756
rect 150308 79716 150342 79756
rect 150308 79704 150314 79716
rect 150434 79704 150440 79756
rect 150492 79716 150526 79756
rect 150492 79704 150498 79716
rect 149848 79580 149974 79608
rect 149848 79568 149854 79580
rect 149698 79540 149704 79552
rect 149164 79512 149704 79540
rect 149698 79500 149704 79512
rect 149756 79500 149762 79552
rect 150590 79540 150618 79988
rect 151326 79960 151354 79988
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 151124 79908 151130 79960
rect 151182 79908 151188 79960
rect 151308 79908 151314 79960
rect 151366 79908 151372 79960
rect 151400 79908 151406 79960
rect 151458 79908 151464 79960
rect 151584 79908 151590 79960
rect 151642 79948 151648 79960
rect 151642 79908 151676 79948
rect 150756 79840 150762 79892
rect 150814 79840 150820 79892
rect 150774 79620 150802 79840
rect 151050 79620 151078 79908
rect 151142 79812 151170 79908
rect 151262 79812 151268 79824
rect 151142 79784 151268 79812
rect 151262 79772 151268 79784
rect 151320 79772 151326 79824
rect 151418 79676 151446 79908
rect 151538 79676 151544 79688
rect 151418 79648 151544 79676
rect 151538 79636 151544 79648
rect 151596 79636 151602 79688
rect 150774 79580 150808 79620
rect 150802 79568 150808 79580
rect 150860 79568 150866 79620
rect 151050 79580 151084 79620
rect 151078 79568 151084 79580
rect 151136 79568 151142 79620
rect 151648 79552 151676 79908
rect 151832 79552 151860 80056
rect 152890 79960 152918 80056
rect 159882 79960 159910 80600
rect 169634 80560 169662 80600
rect 188338 80588 188344 80640
rect 188396 80628 188402 80640
rect 189902 80628 189908 80640
rect 188396 80600 189908 80628
rect 188396 80588 188402 80600
rect 189902 80588 189908 80600
rect 189960 80588 189966 80640
rect 161446 80532 169662 80560
rect 169726 80532 175366 80560
rect 160204 79988 161106 80016
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152780 79908 152786 79960
rect 152838 79908 152844 79960
rect 152872 79908 152878 79960
rect 152930 79908 152936 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 154160 79908 154166 79960
rect 154218 79908 154224 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 154896 79908 154902 79960
rect 154954 79908 154960 79960
rect 154988 79908 154994 79960
rect 155046 79908 155052 79960
rect 155080 79908 155086 79960
rect 155138 79908 155144 79960
rect 155264 79908 155270 79960
rect 155322 79908 155328 79960
rect 155356 79908 155362 79960
rect 155414 79908 155420 79960
rect 155632 79908 155638 79960
rect 155690 79908 155696 79960
rect 155724 79908 155730 79960
rect 155782 79908 155788 79960
rect 155816 79908 155822 79960
rect 155874 79908 155880 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156000 79908 156006 79960
rect 156058 79908 156064 79960
rect 156092 79908 156098 79960
rect 156150 79908 156156 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156644 79908 156650 79960
rect 156702 79908 156708 79960
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157288 79908 157294 79960
rect 157346 79908 157352 79960
rect 158116 79908 158122 79960
rect 158174 79908 158180 79960
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 158576 79908 158582 79960
rect 158634 79908 158640 79960
rect 158668 79908 158674 79960
rect 158726 79908 158732 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 159404 79908 159410 79960
rect 159462 79908 159468 79960
rect 159680 79908 159686 79960
rect 159738 79908 159744 79960
rect 159864 79908 159870 79960
rect 159922 79908 159928 79960
rect 159956 79908 159962 79960
rect 160014 79908 160020 79960
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 151952 79880 151958 79892
rect 151924 79840 151958 79880
rect 152010 79840 152016 79892
rect 152044 79840 152050 79892
rect 152102 79880 152108 79892
rect 152102 79840 152136 79880
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 150710 79540 150716 79552
rect 150590 79512 150716 79540
rect 150710 79500 150716 79512
rect 150768 79500 150774 79552
rect 151630 79500 151636 79552
rect 151688 79500 151694 79552
rect 151814 79500 151820 79552
rect 151872 79500 151878 79552
rect 151924 79472 151952 79840
rect 141068 79444 141188 79472
rect 141160 79404 141188 79444
rect 141344 79444 151952 79472
rect 141344 79404 141372 79444
rect 134076 79376 141004 79404
rect 141160 79376 141372 79404
rect 133840 79364 133846 79376
rect 3510 79296 3516 79348
rect 3568 79336 3574 79348
rect 140774 79336 140780 79348
rect 3568 79308 140780 79336
rect 3568 79296 3574 79308
rect 140774 79296 140780 79308
rect 140832 79296 140838 79348
rect 112254 79228 112260 79280
rect 112312 79268 112318 79280
rect 134426 79268 134432 79280
rect 112312 79240 134432 79268
rect 112312 79228 112318 79240
rect 134426 79228 134432 79240
rect 134484 79228 134490 79280
rect 139486 79228 139492 79280
rect 139544 79268 139550 79280
rect 140498 79268 140504 79280
rect 139544 79240 140504 79268
rect 139544 79228 139550 79240
rect 140498 79228 140504 79240
rect 140556 79228 140562 79280
rect 140976 79268 141004 79376
rect 141418 79364 141424 79416
rect 141476 79404 141482 79416
rect 151170 79404 151176 79416
rect 141476 79376 151176 79404
rect 141476 79364 141482 79376
rect 151170 79364 151176 79376
rect 151228 79364 151234 79416
rect 151906 79364 151912 79416
rect 151964 79404 151970 79416
rect 152108 79404 152136 79840
rect 152246 79756 152274 79840
rect 152182 79704 152188 79756
rect 152240 79716 152274 79756
rect 152240 79704 152246 79716
rect 152430 79676 152458 79908
rect 152688 79880 152694 79892
rect 152660 79840 152694 79880
rect 152746 79840 152752 79892
rect 152798 79880 152826 79908
rect 152964 79880 152970 79892
rect 152798 79852 152872 79880
rect 152660 79756 152688 79840
rect 152642 79704 152648 79756
rect 152700 79704 152706 79756
rect 152844 79688 152872 79852
rect 152936 79840 152970 79880
rect 153022 79840 153028 79892
rect 152936 79688 152964 79840
rect 153010 79704 153016 79756
rect 153068 79744 153074 79756
rect 153166 79744 153194 79908
rect 153240 79840 153246 79892
rect 153298 79840 153304 79892
rect 153068 79716 153194 79744
rect 153068 79704 153074 79716
rect 152430 79648 152780 79676
rect 152642 79432 152648 79484
rect 152700 79472 152706 79484
rect 152752 79472 152780 79648
rect 152826 79636 152832 79688
rect 152884 79636 152890 79688
rect 152918 79636 152924 79688
rect 152976 79636 152982 79688
rect 153102 79636 153108 79688
rect 153160 79676 153166 79688
rect 153258 79676 153286 79840
rect 153442 79756 153470 79908
rect 153792 79840 153798 79892
rect 153850 79840 153856 79892
rect 153976 79880 153982 79892
rect 153948 79840 153982 79880
rect 154034 79840 154040 79892
rect 153442 79716 153476 79756
rect 153470 79704 153476 79716
rect 153528 79704 153534 79756
rect 153810 79688 153838 79840
rect 153948 79756 153976 79840
rect 154178 79812 154206 79908
rect 154040 79784 154206 79812
rect 153930 79704 153936 79756
rect 153988 79704 153994 79756
rect 153378 79676 153384 79688
rect 153160 79636 153194 79676
rect 153258 79648 153384 79676
rect 153378 79636 153384 79648
rect 153436 79636 153442 79688
rect 153746 79636 153752 79688
rect 153804 79648 153838 79688
rect 153804 79636 153810 79648
rect 152700 79444 152780 79472
rect 153166 79472 153194 79636
rect 154040 79608 154068 79784
rect 154114 79704 154120 79756
rect 154172 79744 154178 79756
rect 154270 79744 154298 79908
rect 154172 79716 154298 79744
rect 154172 79704 154178 79716
rect 154638 79688 154666 79908
rect 154804 79880 154810 79892
rect 154776 79840 154810 79880
rect 154862 79840 154868 79892
rect 154776 79688 154804 79840
rect 154914 79756 154942 79908
rect 154850 79704 154856 79756
rect 154908 79716 154942 79756
rect 154908 79704 154914 79716
rect 154574 79636 154580 79688
rect 154632 79648 154666 79688
rect 154632 79636 154638 79648
rect 154758 79636 154764 79688
rect 154816 79636 154822 79688
rect 154666 79608 154672 79620
rect 154040 79580 154672 79608
rect 154666 79568 154672 79580
rect 154724 79568 154730 79620
rect 153930 79472 153936 79484
rect 153166 79444 153936 79472
rect 152700 79432 152706 79444
rect 153930 79432 153936 79444
rect 153988 79432 153994 79484
rect 151964 79376 152136 79404
rect 151964 79364 151970 79376
rect 154298 79364 154304 79416
rect 154356 79404 154362 79416
rect 155006 79404 155034 79908
rect 155098 79688 155126 79908
rect 155098 79648 155132 79688
rect 155126 79636 155132 79648
rect 155184 79636 155190 79688
rect 155282 79540 155310 79908
rect 155374 79620 155402 79908
rect 155650 79880 155678 79908
rect 155604 79852 155678 79880
rect 155604 79824 155632 79852
rect 155448 79772 155454 79824
rect 155506 79772 155512 79824
rect 155586 79772 155592 79824
rect 155644 79772 155650 79824
rect 155742 79812 155770 79908
rect 155696 79784 155770 79812
rect 155466 79688 155494 79772
rect 155696 79688 155724 79784
rect 155834 79756 155862 79908
rect 155926 79824 155954 79908
rect 155908 79772 155914 79824
rect 155966 79772 155972 79824
rect 155770 79704 155776 79756
rect 155828 79716 155862 79756
rect 155828 79704 155834 79716
rect 155466 79648 155500 79688
rect 155494 79636 155500 79648
rect 155552 79636 155558 79688
rect 155678 79636 155684 79688
rect 155736 79636 155742 79688
rect 155862 79636 155868 79688
rect 155920 79676 155926 79688
rect 156018 79676 156046 79908
rect 156110 79756 156138 79908
rect 156202 79812 156230 79908
rect 156202 79784 156276 79812
rect 156110 79716 156144 79756
rect 156138 79704 156144 79716
rect 156196 79704 156202 79756
rect 155920 79648 156046 79676
rect 155920 79636 155926 79648
rect 155374 79580 155408 79620
rect 155402 79568 155408 79580
rect 155460 79568 155466 79620
rect 156248 79608 156276 79784
rect 156386 79688 156414 79908
rect 156460 79772 156466 79824
rect 156518 79772 156524 79824
rect 156322 79636 156328 79688
rect 156380 79648 156414 79688
rect 156478 79688 156506 79772
rect 156478 79648 156512 79688
rect 156380 79636 156386 79648
rect 156506 79636 156512 79648
rect 156564 79636 156570 79688
rect 156414 79608 156420 79620
rect 156248 79580 156420 79608
rect 156414 79568 156420 79580
rect 156472 79568 156478 79620
rect 156662 79552 156690 79908
rect 155954 79540 155960 79552
rect 155282 79512 155960 79540
rect 155954 79500 155960 79512
rect 156012 79500 156018 79552
rect 156598 79500 156604 79552
rect 156656 79512 156690 79552
rect 156656 79500 156662 79512
rect 156938 79472 156966 79908
rect 157214 79880 157242 79908
rect 157168 79852 157242 79880
rect 157168 79540 157196 79852
rect 157306 79756 157334 79908
rect 157472 79840 157478 79892
rect 157530 79840 157536 79892
rect 157932 79840 157938 79892
rect 157990 79840 157996 79892
rect 157242 79704 157248 79756
rect 157300 79716 157334 79756
rect 157300 79704 157306 79716
rect 157490 79608 157518 79840
rect 157610 79704 157616 79756
rect 157668 79704 157674 79756
rect 157950 79744 157978 79840
rect 158134 79824 158162 79908
rect 158134 79784 158168 79824
rect 158162 79772 158168 79784
rect 158220 79772 158226 79824
rect 157950 79716 158116 79744
rect 157628 79676 157656 79704
rect 157978 79676 157984 79688
rect 157628 79648 157984 79676
rect 157978 79636 157984 79648
rect 158036 79636 158042 79688
rect 157610 79608 157616 79620
rect 157490 79580 157616 79608
rect 157610 79568 157616 79580
rect 157668 79568 157674 79620
rect 157702 79540 157708 79552
rect 157168 79512 157708 79540
rect 157702 79500 157708 79512
rect 157760 79500 157766 79552
rect 157334 79472 157340 79484
rect 156938 79444 157340 79472
rect 157334 79432 157340 79444
rect 157392 79432 157398 79484
rect 154356 79376 155034 79404
rect 154356 79364 154362 79376
rect 141234 79296 141240 79348
rect 141292 79336 141298 79348
rect 152458 79336 152464 79348
rect 141292 79308 152464 79336
rect 141292 79296 141298 79308
rect 152458 79296 152464 79308
rect 152516 79296 152522 79348
rect 157426 79296 157432 79348
rect 157484 79336 157490 79348
rect 158088 79336 158116 79716
rect 158502 79620 158530 79908
rect 158438 79568 158444 79620
rect 158496 79580 158530 79620
rect 158496 79568 158502 79580
rect 158594 79552 158622 79908
rect 158686 79744 158714 79908
rect 158760 79772 158766 79824
rect 158818 79812 158824 79824
rect 158818 79784 159036 79812
rect 158818 79772 158824 79784
rect 158686 79716 158852 79744
rect 158824 79688 158852 79716
rect 158806 79636 158812 79688
rect 158864 79636 158870 79688
rect 159008 79552 159036 79784
rect 159330 79756 159358 79908
rect 159422 79812 159450 79908
rect 159422 79784 159496 79812
rect 159330 79716 159364 79756
rect 159358 79704 159364 79716
rect 159416 79704 159422 79756
rect 158530 79500 158536 79552
rect 158588 79512 158622 79552
rect 158898 79540 158904 79552
rect 158686 79512 158904 79540
rect 158588 79500 158594 79512
rect 158254 79432 158260 79484
rect 158312 79472 158318 79484
rect 158686 79472 158714 79512
rect 158898 79500 158904 79512
rect 158956 79500 158962 79552
rect 158990 79500 158996 79552
rect 159048 79500 159054 79552
rect 158312 79444 158714 79472
rect 158312 79432 158318 79444
rect 158898 79364 158904 79416
rect 158956 79404 158962 79416
rect 159468 79404 159496 79784
rect 159588 79772 159594 79824
rect 159646 79772 159652 79824
rect 159606 79688 159634 79772
rect 159542 79636 159548 79688
rect 159600 79648 159634 79688
rect 159600 79636 159606 79648
rect 159698 79620 159726 79908
rect 159634 79568 159640 79620
rect 159692 79580 159726 79620
rect 159974 79608 160002 79908
rect 159836 79580 160002 79608
rect 159692 79568 159698 79580
rect 159836 79552 159864 79580
rect 160066 79552 160094 79908
rect 160204 79620 160232 79988
rect 161078 79960 161106 79988
rect 161446 79960 161474 80532
rect 163102 79988 163452 80016
rect 163102 79960 163130 79988
rect 160324 79908 160330 79960
rect 160382 79908 160388 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160508 79908 160514 79960
rect 160566 79908 160572 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160692 79908 160698 79960
rect 160750 79908 160756 79960
rect 160784 79908 160790 79960
rect 160842 79908 160848 79960
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 161060 79908 161066 79960
rect 161118 79908 161124 79960
rect 161428 79908 161434 79960
rect 161486 79908 161492 79960
rect 161612 79908 161618 79960
rect 161670 79908 161676 79960
rect 161704 79908 161710 79960
rect 161762 79908 161768 79960
rect 161796 79908 161802 79960
rect 161854 79908 161860 79960
rect 161980 79908 161986 79960
rect 162038 79948 162044 79960
rect 162038 79908 162072 79948
rect 162440 79908 162446 79960
rect 162498 79908 162504 79960
rect 162532 79908 162538 79960
rect 162590 79948 162596 79960
rect 162590 79908 162624 79948
rect 162808 79908 162814 79960
rect 162866 79948 162872 79960
rect 162866 79908 162900 79948
rect 162992 79908 162998 79960
rect 163050 79908 163056 79960
rect 163084 79908 163090 79960
rect 163142 79908 163148 79960
rect 163268 79908 163274 79960
rect 163326 79908 163332 79960
rect 160186 79568 160192 79620
rect 160244 79568 160250 79620
rect 159818 79500 159824 79552
rect 159876 79500 159882 79552
rect 160002 79500 160008 79552
rect 160060 79512 160094 79552
rect 160060 79500 160066 79512
rect 158956 79376 159496 79404
rect 160342 79404 160370 79908
rect 160434 79688 160462 79908
rect 160526 79824 160554 79908
rect 160508 79772 160514 79824
rect 160566 79772 160572 79824
rect 160434 79648 160468 79688
rect 160462 79636 160468 79648
rect 160520 79636 160526 79688
rect 160618 79620 160646 79908
rect 160710 79676 160738 79908
rect 160802 79744 160830 79908
rect 160894 79812 160922 79908
rect 160894 79784 161244 79812
rect 161106 79744 161112 79756
rect 160802 79716 161112 79744
rect 161106 79704 161112 79716
rect 161164 79704 161170 79756
rect 160830 79676 160836 79688
rect 160710 79648 160836 79676
rect 160830 79636 160836 79648
rect 160888 79636 160894 79688
rect 161216 79620 161244 79784
rect 161630 79620 161658 79908
rect 161722 79756 161750 79908
rect 161814 79812 161842 79908
rect 161888 79840 161894 79892
rect 161946 79880 161952 79892
rect 161946 79840 161980 79880
rect 161814 79784 161888 79812
rect 161860 79756 161888 79784
rect 161722 79716 161756 79756
rect 161750 79704 161756 79716
rect 161808 79704 161814 79756
rect 161842 79704 161848 79756
rect 161900 79704 161906 79756
rect 160618 79580 160652 79620
rect 160646 79568 160652 79580
rect 160704 79568 160710 79620
rect 161198 79568 161204 79620
rect 161256 79568 161262 79620
rect 161630 79580 161664 79620
rect 161658 79568 161664 79580
rect 161716 79568 161722 79620
rect 161566 79500 161572 79552
rect 161624 79540 161630 79552
rect 161952 79540 161980 79840
rect 162044 79552 162072 79908
rect 162458 79880 162486 79908
rect 162458 79852 162532 79880
rect 162504 79756 162532 79852
rect 162486 79704 162492 79756
rect 162544 79704 162550 79756
rect 162596 79608 162624 79908
rect 162716 79812 162722 79824
rect 162688 79772 162722 79812
rect 162774 79772 162780 79824
rect 162688 79688 162716 79772
rect 162670 79636 162676 79688
rect 162728 79636 162734 79688
rect 162762 79608 162768 79620
rect 162596 79580 162768 79608
rect 162762 79568 162768 79580
rect 162820 79568 162826 79620
rect 161624 79512 161980 79540
rect 161624 79500 161630 79512
rect 162026 79500 162032 79552
rect 162084 79500 162090 79552
rect 162872 79472 162900 79908
rect 163010 79824 163038 79908
rect 163010 79784 163044 79824
rect 163038 79772 163044 79784
rect 163096 79772 163102 79824
rect 163286 79552 163314 79908
rect 163424 79688 163452 79988
rect 168898 79988 169662 80016
rect 168898 79960 168926 79988
rect 163636 79908 163642 79960
rect 163694 79908 163700 79960
rect 163820 79908 163826 79960
rect 163878 79908 163884 79960
rect 164096 79908 164102 79960
rect 164154 79908 164160 79960
rect 164556 79908 164562 79960
rect 164614 79908 164620 79960
rect 164648 79908 164654 79960
rect 164706 79908 164712 79960
rect 164740 79908 164746 79960
rect 164798 79908 164804 79960
rect 164924 79908 164930 79960
rect 164982 79908 164988 79960
rect 165016 79908 165022 79960
rect 165074 79908 165080 79960
rect 165200 79948 165206 79960
rect 165172 79908 165206 79948
rect 165258 79908 165264 79960
rect 165384 79948 165390 79960
rect 165356 79908 165390 79948
rect 165442 79908 165448 79960
rect 165660 79908 165666 79960
rect 165718 79908 165724 79960
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 166396 79948 166402 79960
rect 166230 79920 166402 79948
rect 163654 79880 163682 79908
rect 163608 79852 163682 79880
rect 163406 79636 163412 79688
rect 163464 79636 163470 79688
rect 163608 79620 163636 79852
rect 163728 79840 163734 79892
rect 163786 79840 163792 79892
rect 163746 79688 163774 79840
rect 163838 79824 163866 79908
rect 163838 79784 163872 79824
rect 163866 79772 163872 79784
rect 163924 79772 163930 79824
rect 164114 79688 164142 79908
rect 164372 79840 164378 79892
rect 164430 79840 164436 79892
rect 164188 79772 164194 79824
rect 164246 79772 164252 79824
rect 163682 79636 163688 79688
rect 163740 79648 163774 79688
rect 163740 79636 163746 79648
rect 164050 79636 164056 79688
rect 164108 79648 164142 79688
rect 164206 79688 164234 79772
rect 164206 79648 164240 79688
rect 164108 79636 164114 79648
rect 164234 79636 164240 79648
rect 164292 79636 164298 79688
rect 164390 79620 164418 79840
rect 164574 79756 164602 79908
rect 164510 79704 164516 79756
rect 164568 79716 164602 79756
rect 164568 79704 164574 79716
rect 164666 79620 164694 79908
rect 163590 79568 163596 79620
rect 163648 79568 163654 79620
rect 164390 79580 164424 79620
rect 164418 79568 164424 79580
rect 164476 79568 164482 79620
rect 164602 79568 164608 79620
rect 164660 79580 164694 79620
rect 164660 79568 164666 79580
rect 164758 79552 164786 79908
rect 164942 79880 164970 79908
rect 164896 79852 164970 79880
rect 164896 79688 164924 79852
rect 165034 79756 165062 79908
rect 165172 79756 165200 79908
rect 165356 79824 165384 79908
rect 165568 79880 165574 79892
rect 165448 79852 165574 79880
rect 165338 79772 165344 79824
rect 165396 79772 165402 79824
rect 164970 79704 164976 79756
rect 165028 79716 165062 79756
rect 165028 79704 165034 79716
rect 165154 79704 165160 79756
rect 165212 79704 165218 79756
rect 164878 79636 164884 79688
rect 164936 79636 164942 79688
rect 165448 79620 165476 79852
rect 165568 79840 165574 79852
rect 165626 79840 165632 79892
rect 165678 79756 165706 79908
rect 165614 79704 165620 79756
rect 165672 79716 165706 79756
rect 165770 79756 165798 79908
rect 165936 79880 165942 79892
rect 165908 79840 165942 79880
rect 165994 79840 166000 79892
rect 165770 79716 165804 79756
rect 165672 79704 165678 79716
rect 165798 79704 165804 79716
rect 165856 79704 165862 79756
rect 165908 79688 165936 79840
rect 166120 79772 166126 79824
rect 166178 79772 166184 79824
rect 166138 79688 166166 79772
rect 165890 79636 165896 79688
rect 165948 79636 165954 79688
rect 166074 79636 166080 79688
rect 166132 79648 166166 79688
rect 166132 79636 166138 79648
rect 165430 79568 165436 79620
rect 165488 79568 165494 79620
rect 166230 79608 166258 79920
rect 166396 79908 166402 79920
rect 166454 79908 166460 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166764 79908 166770 79960
rect 166822 79908 166828 79960
rect 167132 79908 167138 79960
rect 167190 79908 167196 79960
rect 167224 79908 167230 79960
rect 167282 79908 167288 79960
rect 167500 79948 167506 79960
rect 167472 79908 167506 79948
rect 167558 79908 167564 79960
rect 167684 79908 167690 79960
rect 167742 79908 167748 79960
rect 167776 79908 167782 79960
rect 167834 79908 167840 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168788 79908 168794 79960
rect 168846 79908 168852 79960
rect 168880 79908 168886 79960
rect 168938 79908 168944 79960
rect 168972 79908 168978 79960
rect 169030 79908 169036 79960
rect 169064 79908 169070 79960
rect 169122 79908 169128 79960
rect 169340 79908 169346 79960
rect 169398 79908 169404 79960
rect 166304 79772 166310 79824
rect 166362 79772 166368 79824
rect 166322 79688 166350 79772
rect 166506 79688 166534 79908
rect 166690 79756 166718 79908
rect 166626 79704 166632 79756
rect 166684 79716 166718 79756
rect 166684 79704 166690 79716
rect 166322 79648 166356 79688
rect 166350 79636 166356 79648
rect 166408 79636 166414 79688
rect 166442 79636 166448 79688
rect 166500 79648 166534 79688
rect 166500 79636 166506 79648
rect 166534 79608 166540 79620
rect 166230 79580 166540 79608
rect 166534 79568 166540 79580
rect 166592 79568 166598 79620
rect 166782 79608 166810 79908
rect 167150 79620 167178 79908
rect 167242 79812 167270 79908
rect 167316 79840 167322 79892
rect 167374 79880 167380 79892
rect 167374 79840 167408 79880
rect 167242 79784 167316 79812
rect 167288 79756 167316 79784
rect 167270 79704 167276 79756
rect 167328 79704 167334 79756
rect 167380 79620 167408 79840
rect 167472 79688 167500 79908
rect 167592 79840 167598 79892
rect 167650 79840 167656 79892
rect 167454 79636 167460 79688
rect 167512 79636 167518 79688
rect 167610 79620 167638 79840
rect 166994 79608 167000 79620
rect 166782 79580 167000 79608
rect 166994 79568 167000 79580
rect 167052 79568 167058 79620
rect 167150 79580 167184 79620
rect 167178 79568 167184 79580
rect 167236 79568 167242 79620
rect 167362 79568 167368 79620
rect 167420 79568 167426 79620
rect 167546 79568 167552 79620
rect 167604 79580 167638 79620
rect 167604 79568 167610 79580
rect 163286 79512 163320 79552
rect 163314 79500 163320 79512
rect 163372 79500 163378 79552
rect 164694 79500 164700 79552
rect 164752 79512 164786 79552
rect 167702 79540 167730 79908
rect 167794 79620 167822 79908
rect 168438 79688 168466 79908
rect 168512 79840 168518 79892
rect 168570 79880 168576 79892
rect 168570 79840 168604 79880
rect 168438 79648 168472 79688
rect 168466 79636 168472 79648
rect 168524 79636 168530 79688
rect 168576 79620 168604 79840
rect 168806 79756 168834 79908
rect 168990 79824 169018 79908
rect 168926 79772 168932 79824
rect 168984 79784 169018 79824
rect 168984 79772 168990 79784
rect 168806 79716 168840 79756
rect 168834 79704 168840 79716
rect 168892 79704 168898 79756
rect 169082 79620 169110 79908
rect 167794 79580 167828 79620
rect 167822 79568 167828 79580
rect 167880 79568 167886 79620
rect 168558 79568 168564 79620
rect 168616 79568 168622 79620
rect 169018 79568 169024 79620
rect 169076 79580 169110 79620
rect 169358 79620 169386 79908
rect 169634 79824 169662 79988
rect 169726 79960 169754 80532
rect 175338 80492 175366 80532
rect 186958 80520 186964 80572
rect 187016 80560 187022 80572
rect 192662 80560 192668 80572
rect 187016 80532 192668 80560
rect 187016 80520 187022 80532
rect 192662 80520 192668 80532
rect 192720 80520 192726 80572
rect 179598 80492 179604 80504
rect 175016 80464 175228 80492
rect 175338 80464 179604 80492
rect 175016 80424 175044 80464
rect 173038 80396 175044 80424
rect 175200 80424 175228 80464
rect 179598 80452 179604 80464
rect 179656 80452 179662 80504
rect 187050 80452 187056 80504
rect 187108 80492 187114 80504
rect 191098 80492 191104 80504
rect 187108 80464 191104 80492
rect 187108 80452 187114 80464
rect 191098 80452 191104 80464
rect 191156 80452 191162 80504
rect 178126 80424 178132 80436
rect 175200 80396 178132 80424
rect 173038 79960 173066 80396
rect 178126 80384 178132 80396
rect 178184 80384 178190 80436
rect 175246 80328 178034 80356
rect 175246 80288 175274 80328
rect 174326 80260 175274 80288
rect 178006 80300 178034 80328
rect 178006 80260 178040 80300
rect 174326 80016 174354 80260
rect 178034 80248 178040 80260
rect 178092 80248 178098 80300
rect 173130 79988 174354 80016
rect 174970 80192 177712 80220
rect 169708 79908 169714 79960
rect 169766 79908 169772 79960
rect 169892 79908 169898 79960
rect 169950 79908 169956 79960
rect 170168 79908 170174 79960
rect 170226 79908 170232 79960
rect 170444 79908 170450 79960
rect 170502 79908 170508 79960
rect 170536 79908 170542 79960
rect 170594 79908 170600 79960
rect 171272 79908 171278 79960
rect 171330 79908 171336 79960
rect 171640 79948 171646 79960
rect 171612 79908 171646 79948
rect 171698 79908 171704 79960
rect 172100 79908 172106 79960
rect 172158 79908 172164 79960
rect 172192 79908 172198 79960
rect 172250 79908 172256 79960
rect 172376 79908 172382 79960
rect 172434 79908 172440 79960
rect 172560 79908 172566 79960
rect 172618 79908 172624 79960
rect 173020 79908 173026 79960
rect 173078 79908 173084 79960
rect 169634 79784 169668 79824
rect 169662 79772 169668 79784
rect 169720 79772 169726 79824
rect 169910 79812 169938 79908
rect 169772 79784 169938 79812
rect 169772 79676 169800 79784
rect 170186 79688 170214 79908
rect 170352 79880 170358 79892
rect 170324 79840 170358 79880
rect 170410 79840 170416 79892
rect 170324 79756 170352 79840
rect 170462 79756 170490 79908
rect 170306 79704 170312 79756
rect 170364 79704 170370 79756
rect 170398 79704 170404 79756
rect 170456 79716 170490 79756
rect 170456 79704 170462 79716
rect 170554 79688 170582 79908
rect 170996 79840 171002 79892
rect 171054 79840 171060 79892
rect 171180 79840 171186 79892
rect 171238 79840 171244 79892
rect 171014 79688 171042 79840
rect 170030 79676 170036 79688
rect 169772 79648 170036 79676
rect 170030 79636 170036 79648
rect 170088 79636 170094 79688
rect 170122 79636 170128 79688
rect 170180 79648 170214 79688
rect 170180 79636 170186 79648
rect 170490 79636 170496 79688
rect 170548 79648 170582 79688
rect 170548 79636 170554 79648
rect 170950 79636 170956 79688
rect 171008 79648 171042 79688
rect 171008 79636 171014 79648
rect 169358 79580 169392 79620
rect 169076 79568 169082 79580
rect 169386 79568 169392 79580
rect 169444 79568 169450 79620
rect 167914 79540 167920 79552
rect 167702 79512 167920 79540
rect 164752 79500 164758 79512
rect 167914 79500 167920 79512
rect 167972 79500 167978 79552
rect 165614 79472 165620 79484
rect 162872 79444 165620 79472
rect 165614 79432 165620 79444
rect 165672 79432 165678 79484
rect 162578 79404 162584 79416
rect 160342 79376 162584 79404
rect 158956 79364 158962 79376
rect 162578 79364 162584 79376
rect 162636 79364 162642 79416
rect 162826 79376 165614 79404
rect 157484 79308 158116 79336
rect 157484 79296 157490 79308
rect 141418 79268 141424 79280
rect 140976 79240 141424 79268
rect 141418 79228 141424 79240
rect 141476 79228 141482 79280
rect 145282 79228 145288 79280
rect 145340 79268 145346 79280
rect 145558 79268 145564 79280
rect 145340 79240 145564 79268
rect 145340 79228 145346 79240
rect 145558 79228 145564 79240
rect 145616 79228 145622 79280
rect 162826 79268 162854 79376
rect 165586 79336 165614 79376
rect 166534 79364 166540 79416
rect 166592 79404 166598 79416
rect 168282 79404 168288 79416
rect 166592 79376 168288 79404
rect 166592 79364 166598 79376
rect 168282 79364 168288 79376
rect 168340 79364 168346 79416
rect 171198 79404 171226 79840
rect 171290 79608 171318 79908
rect 171612 79688 171640 79908
rect 171824 79840 171830 79892
rect 171882 79840 171888 79892
rect 171594 79636 171600 79688
rect 171652 79636 171658 79688
rect 171842 79676 171870 79840
rect 171962 79676 171968 79688
rect 171842 79648 171968 79676
rect 171962 79636 171968 79648
rect 172020 79636 172026 79688
rect 172118 79676 172146 79908
rect 172210 79756 172238 79908
rect 172394 79824 172422 79908
rect 172578 79880 172606 79908
rect 173130 79880 173158 79988
rect 174970 79960 174998 80192
rect 177684 80084 177712 80192
rect 177758 80180 177764 80232
rect 177816 80220 177822 80232
rect 178954 80220 178960 80232
rect 177816 80192 178960 80220
rect 177816 80180 177822 80192
rect 178954 80180 178960 80192
rect 179012 80180 179018 80232
rect 179230 80084 179236 80096
rect 177684 80056 179236 80084
rect 179230 80044 179236 80056
rect 179288 80044 179294 80096
rect 203794 80044 203800 80096
rect 203852 80084 203858 80096
rect 204714 80084 204720 80096
rect 203852 80056 204720 80084
rect 203852 80044 203858 80056
rect 204714 80044 204720 80056
rect 204772 80044 204778 80096
rect 182818 80016 182824 80028
rect 176166 79988 182824 80016
rect 176166 79960 176194 79988
rect 182818 79976 182824 79988
rect 182876 79976 182882 80028
rect 183922 79976 183928 80028
rect 183980 80016 183986 80028
rect 190822 80016 190828 80028
rect 183980 79988 190828 80016
rect 183980 79976 183986 79988
rect 190822 79976 190828 79988
rect 190880 79976 190886 80028
rect 202322 79976 202328 80028
rect 202380 80016 202386 80028
rect 202782 80016 202788 80028
rect 202380 79988 202788 80016
rect 202380 79976 202386 79988
rect 202782 79976 202788 79988
rect 202840 80016 202846 80028
rect 580166 80016 580172 80028
rect 202840 79988 580172 80016
rect 202840 79976 202846 79988
rect 580166 79976 580172 79988
rect 580224 79976 580230 80028
rect 173756 79908 173762 79960
rect 173814 79948 173820 79960
rect 173814 79920 173940 79948
rect 173814 79908 173820 79920
rect 172578 79852 172652 79880
rect 172624 79824 172652 79852
rect 172716 79852 173158 79880
rect 172394 79784 172428 79824
rect 172422 79772 172428 79784
rect 172480 79772 172486 79824
rect 172606 79772 172612 79824
rect 172664 79772 172670 79824
rect 172210 79716 172244 79756
rect 172238 79704 172244 79716
rect 172296 79704 172302 79756
rect 172330 79676 172336 79688
rect 172118 79648 172336 79676
rect 172330 79636 172336 79648
rect 172388 79636 172394 79688
rect 171778 79608 171784 79620
rect 171290 79580 171784 79608
rect 171778 79568 171784 79580
rect 171836 79568 171842 79620
rect 172716 79540 172744 79852
rect 173204 79840 173210 79892
rect 173262 79840 173268 79892
rect 173572 79840 173578 79892
rect 173630 79840 173636 79892
rect 173222 79676 173250 79840
rect 173388 79772 173394 79824
rect 173446 79772 173452 79824
rect 173590 79812 173618 79840
rect 173590 79784 173664 79812
rect 171520 79512 172744 79540
rect 173176 79648 173250 79676
rect 173406 79688 173434 79772
rect 173406 79648 173440 79688
rect 173176 79540 173204 79648
rect 173434 79636 173440 79648
rect 173492 79636 173498 79688
rect 173636 79620 173664 79784
rect 173912 79688 173940 79920
rect 174860 79908 174866 79960
rect 174918 79908 174924 79960
rect 174952 79908 174958 79960
rect 175010 79908 175016 79960
rect 175412 79908 175418 79960
rect 175470 79908 175476 79960
rect 175872 79908 175878 79960
rect 175930 79948 175936 79960
rect 175930 79920 176056 79948
rect 175930 79908 175936 79920
rect 174032 79880 174038 79892
rect 174004 79840 174038 79880
rect 174090 79840 174096 79892
rect 174124 79840 174130 79892
rect 174182 79880 174188 79892
rect 174878 79880 174906 79908
rect 175136 79880 175142 79892
rect 174182 79852 174814 79880
rect 174878 79852 174952 79880
rect 174182 79840 174188 79852
rect 173894 79636 173900 79688
rect 173952 79636 173958 79688
rect 174004 79620 174032 79840
rect 174492 79772 174498 79824
rect 174550 79772 174556 79824
rect 174584 79772 174590 79824
rect 174642 79772 174648 79824
rect 174510 79620 174538 79772
rect 174602 79676 174630 79772
rect 174786 79744 174814 79852
rect 174924 79824 174952 79852
rect 175016 79852 175142 79880
rect 174906 79772 174912 79824
rect 174964 79772 174970 79824
rect 174786 79716 174952 79744
rect 174814 79676 174820 79688
rect 174602 79648 174820 79676
rect 174814 79636 174820 79648
rect 174872 79636 174878 79688
rect 173250 79568 173256 79620
rect 173308 79608 173314 79620
rect 173526 79608 173532 79620
rect 173308 79580 173532 79608
rect 173308 79568 173314 79580
rect 173526 79568 173532 79580
rect 173584 79568 173590 79620
rect 173618 79568 173624 79620
rect 173676 79568 173682 79620
rect 173986 79568 173992 79620
rect 174044 79568 174050 79620
rect 174510 79580 174544 79620
rect 174538 79568 174544 79580
rect 174596 79568 174602 79620
rect 174924 79608 174952 79716
rect 175016 79688 175044 79852
rect 175136 79840 175142 79852
rect 175194 79840 175200 79892
rect 175320 79880 175326 79892
rect 175292 79840 175326 79880
rect 175378 79840 175384 79892
rect 175292 79688 175320 79840
rect 175430 79756 175458 79908
rect 175780 79840 175786 79892
rect 175838 79880 175844 79892
rect 175838 79840 175872 79880
rect 175504 79772 175510 79824
rect 175562 79772 175568 79824
rect 175596 79772 175602 79824
rect 175654 79772 175660 79824
rect 175366 79704 175372 79756
rect 175424 79716 175458 79756
rect 175424 79704 175430 79716
rect 175522 79688 175550 79772
rect 174998 79636 175004 79688
rect 175056 79636 175062 79688
rect 175274 79636 175280 79688
rect 175332 79636 175338 79688
rect 175458 79636 175464 79688
rect 175516 79648 175550 79688
rect 175614 79688 175642 79772
rect 175844 79756 175872 79840
rect 175826 79704 175832 79756
rect 175884 79704 175890 79756
rect 176028 79688 176056 79920
rect 176148 79908 176154 79960
rect 176206 79908 176212 79960
rect 176240 79908 176246 79960
rect 176298 79908 176304 79960
rect 176424 79908 176430 79960
rect 176482 79948 176488 79960
rect 177850 79948 177856 79960
rect 176482 79920 177856 79948
rect 176482 79908 176488 79920
rect 177850 79908 177856 79920
rect 177908 79908 177914 79960
rect 185578 79908 185584 79960
rect 185636 79948 185642 79960
rect 214282 79948 214288 79960
rect 185636 79920 214288 79948
rect 185636 79908 185642 79920
rect 214282 79908 214288 79920
rect 214340 79908 214346 79960
rect 176258 79824 176286 79908
rect 176700 79840 176706 79892
rect 176758 79840 176764 79892
rect 176792 79840 176798 79892
rect 176850 79840 176856 79892
rect 176976 79840 176982 79892
rect 177034 79840 177040 79892
rect 177068 79840 177074 79892
rect 177126 79840 177132 79892
rect 177160 79840 177166 79892
rect 177218 79880 177224 79892
rect 177758 79880 177764 79892
rect 177218 79852 177764 79880
rect 177218 79840 177224 79852
rect 177758 79840 177764 79852
rect 177816 79840 177822 79892
rect 179046 79880 179052 79892
rect 178006 79852 179052 79880
rect 176194 79772 176200 79824
rect 176252 79784 176286 79824
rect 176252 79772 176258 79784
rect 176718 79744 176746 79840
rect 176580 79716 176746 79744
rect 175614 79648 175648 79688
rect 175516 79636 175522 79648
rect 175642 79636 175648 79648
rect 175700 79636 175706 79688
rect 176010 79636 176016 79688
rect 176068 79636 176074 79688
rect 176286 79608 176292 79620
rect 174924 79580 176292 79608
rect 176286 79568 176292 79580
rect 176344 79568 176350 79620
rect 175918 79540 175924 79552
rect 173176 79512 175924 79540
rect 171410 79404 171416 79416
rect 171198 79376 171416 79404
rect 171410 79364 171416 79376
rect 171468 79364 171474 79416
rect 171520 79336 171548 79512
rect 175918 79500 175924 79512
rect 175976 79500 175982 79552
rect 176580 79540 176608 79716
rect 176654 79568 176660 79620
rect 176712 79608 176718 79620
rect 176810 79608 176838 79840
rect 176712 79580 176838 79608
rect 176712 79568 176718 79580
rect 176994 79552 177022 79840
rect 177086 79812 177114 79840
rect 178006 79812 178034 79852
rect 179046 79840 179052 79852
rect 179104 79840 179110 79892
rect 177086 79784 178034 79812
rect 178034 79704 178040 79756
rect 178092 79744 178098 79756
rect 580626 79744 580632 79756
rect 178092 79716 580632 79744
rect 178092 79704 178098 79716
rect 580626 79704 580632 79716
rect 580684 79704 580690 79756
rect 177114 79568 177120 79620
rect 177172 79608 177178 79620
rect 179782 79608 179788 79620
rect 177172 79580 179788 79608
rect 177172 79568 177178 79580
rect 179782 79568 179788 79580
rect 179840 79568 179846 79620
rect 176838 79540 176844 79552
rect 176580 79512 176844 79540
rect 176838 79500 176844 79512
rect 176896 79500 176902 79552
rect 176994 79512 177028 79552
rect 177022 79500 177028 79512
rect 177080 79500 177086 79552
rect 177390 79500 177396 79552
rect 177448 79540 177454 79552
rect 209130 79540 209136 79552
rect 177448 79512 209136 79540
rect 177448 79500 177454 79512
rect 209130 79500 209136 79512
rect 209188 79500 209194 79552
rect 172054 79432 172060 79484
rect 172112 79472 172118 79484
rect 172698 79472 172704 79484
rect 172112 79444 172704 79472
rect 172112 79432 172118 79444
rect 172698 79432 172704 79444
rect 172756 79432 172762 79484
rect 173526 79432 173532 79484
rect 173584 79472 173590 79484
rect 189166 79472 189172 79484
rect 173584 79444 189172 79472
rect 173584 79432 173590 79444
rect 189166 79432 189172 79444
rect 189224 79432 189230 79484
rect 201862 79404 201868 79416
rect 165586 79308 171548 79336
rect 171612 79376 201868 79404
rect 152936 79240 162854 79268
rect 119430 79160 119436 79212
rect 119488 79200 119494 79212
rect 150342 79200 150348 79212
rect 119488 79172 150348 79200
rect 119488 79160 119494 79172
rect 150342 79160 150348 79172
rect 150400 79160 150406 79212
rect 112438 79092 112444 79144
rect 112496 79132 112502 79144
rect 144914 79132 144920 79144
rect 112496 79104 144920 79132
rect 112496 79092 112502 79104
rect 144914 79092 144920 79104
rect 144972 79092 144978 79144
rect 145282 79092 145288 79144
rect 145340 79132 145346 79144
rect 145742 79132 145748 79144
rect 145340 79104 145748 79132
rect 145340 79092 145346 79104
rect 145742 79092 145748 79104
rect 145800 79092 145806 79144
rect 151170 79092 151176 79144
rect 151228 79132 151234 79144
rect 152936 79132 152964 79240
rect 168098 79228 168104 79280
rect 168156 79268 168162 79280
rect 171612 79268 171640 79376
rect 201862 79364 201868 79376
rect 201920 79364 201926 79416
rect 173526 79336 173532 79348
rect 168156 79240 171640 79268
rect 171842 79308 173532 79336
rect 168156 79228 168162 79240
rect 161474 79160 161480 79212
rect 161532 79200 161538 79212
rect 161532 79172 168374 79200
rect 161532 79160 161538 79172
rect 168346 79132 168374 79172
rect 170674 79160 170680 79212
rect 170732 79200 170738 79212
rect 171042 79200 171048 79212
rect 170732 79172 171048 79200
rect 170732 79160 170738 79172
rect 171042 79160 171048 79172
rect 171100 79160 171106 79212
rect 171842 79132 171870 79308
rect 173526 79296 173532 79308
rect 173584 79296 173590 79348
rect 197998 79336 198004 79348
rect 173866 79308 198004 79336
rect 173866 79268 173894 79308
rect 197998 79296 198004 79308
rect 198056 79296 198062 79348
rect 175366 79268 175372 79280
rect 151228 79104 152964 79132
rect 154546 79104 162854 79132
rect 168346 79104 171870 79132
rect 171934 79240 173894 79268
rect 174832 79240 175372 79268
rect 151228 79092 151234 79104
rect 118050 79024 118056 79076
rect 118108 79064 118114 79076
rect 153010 79064 153016 79076
rect 118108 79036 153016 79064
rect 118108 79024 118114 79036
rect 153010 79024 153016 79036
rect 153068 79024 153074 79076
rect 111242 78956 111248 79008
rect 111300 78996 111306 79008
rect 146110 78996 146116 79008
rect 111300 78968 146116 78996
rect 111300 78956 111306 78968
rect 146110 78956 146116 78968
rect 146168 78956 146174 79008
rect 149054 78956 149060 79008
rect 149112 78996 149118 79008
rect 154546 78996 154574 79104
rect 149112 78968 154574 78996
rect 162826 78996 162854 79104
rect 164234 79024 164240 79076
rect 164292 79064 164298 79076
rect 171934 79064 171962 79240
rect 172146 79160 172152 79212
rect 172204 79200 172210 79212
rect 174832 79200 174860 79240
rect 175366 79228 175372 79240
rect 175424 79228 175430 79280
rect 175550 79228 175556 79280
rect 175608 79268 175614 79280
rect 176286 79268 176292 79280
rect 175608 79240 176292 79268
rect 175608 79228 175614 79240
rect 176286 79228 176292 79240
rect 176344 79228 176350 79280
rect 176470 79228 176476 79280
rect 176528 79268 176534 79280
rect 210418 79268 210424 79280
rect 176528 79240 210424 79268
rect 176528 79228 176534 79240
rect 210418 79228 210424 79240
rect 210476 79228 210482 79280
rect 172204 79172 174860 79200
rect 172204 79160 172210 79172
rect 174906 79160 174912 79212
rect 174964 79200 174970 79212
rect 209222 79200 209228 79212
rect 174964 79172 209228 79200
rect 174964 79160 174970 79172
rect 209222 79160 209228 79172
rect 209280 79160 209286 79212
rect 181346 79132 181352 79144
rect 172118 79104 181352 79132
rect 172118 79064 172146 79104
rect 181346 79092 181352 79104
rect 181404 79092 181410 79144
rect 210602 79132 210608 79144
rect 181548 79104 210608 79132
rect 181438 79064 181444 79076
rect 164292 79036 171962 79064
rect 172026 79036 172146 79064
rect 175246 79036 181444 79064
rect 164292 79024 164298 79036
rect 172026 78996 172054 79036
rect 162826 78968 172054 78996
rect 149112 78956 149118 78968
rect 172882 78956 172888 79008
rect 172940 78996 172946 79008
rect 174078 78996 174084 79008
rect 172940 78968 174084 78996
rect 172940 78956 172946 78968
rect 174078 78956 174084 78968
rect 174136 78956 174142 79008
rect 121914 78888 121920 78940
rect 121972 78928 121978 78940
rect 162670 78928 162676 78940
rect 121972 78900 162676 78928
rect 121972 78888 121978 78900
rect 162670 78888 162676 78900
rect 162728 78888 162734 78940
rect 167914 78888 167920 78940
rect 167972 78928 167978 78940
rect 175246 78928 175274 79036
rect 181438 79024 181444 79036
rect 181496 79024 181502 79076
rect 176746 78956 176752 79008
rect 176804 78996 176810 79008
rect 181548 78996 181576 79104
rect 210602 79092 210608 79104
rect 210660 79092 210666 79144
rect 202782 79064 202788 79076
rect 190426 79036 202788 79064
rect 176804 78968 181576 78996
rect 176804 78956 176810 78968
rect 181622 78956 181628 79008
rect 181680 78996 181686 79008
rect 190426 78996 190454 79036
rect 202782 79024 202788 79036
rect 202840 79024 202846 79076
rect 181680 78968 190454 78996
rect 181680 78956 181686 78968
rect 167972 78900 175274 78928
rect 167972 78888 167978 78900
rect 178126 78888 178132 78940
rect 178184 78928 178190 78940
rect 212718 78928 212724 78940
rect 178184 78900 212724 78928
rect 178184 78888 178190 78900
rect 212718 78888 212724 78900
rect 212776 78888 212782 78940
rect 98822 78820 98828 78872
rect 98880 78860 98886 78872
rect 139578 78860 139584 78872
rect 98880 78832 139584 78860
rect 98880 78820 98886 78832
rect 139578 78820 139584 78832
rect 139636 78820 139642 78872
rect 142338 78820 142344 78872
rect 142396 78860 142402 78872
rect 142982 78860 142988 78872
rect 142396 78832 142988 78860
rect 142396 78820 142402 78832
rect 142982 78820 142988 78832
rect 143040 78820 143046 78872
rect 158346 78820 158352 78872
rect 158404 78860 158410 78872
rect 158714 78860 158720 78872
rect 158404 78832 158720 78860
rect 158404 78820 158410 78832
rect 158714 78820 158720 78832
rect 158772 78820 158778 78872
rect 171134 78820 171140 78872
rect 171192 78860 171198 78872
rect 211522 78860 211528 78872
rect 171192 78832 211528 78860
rect 171192 78820 171198 78832
rect 211522 78820 211528 78832
rect 211580 78820 211586 78872
rect 133322 78752 133328 78804
rect 133380 78792 133386 78804
rect 137002 78792 137008 78804
rect 133380 78764 137008 78792
rect 133380 78752 133386 78764
rect 137002 78752 137008 78764
rect 137060 78752 137066 78804
rect 140498 78752 140504 78804
rect 140556 78792 140562 78804
rect 144638 78792 144644 78804
rect 140556 78764 144644 78792
rect 140556 78752 140562 78764
rect 144638 78752 144644 78764
rect 144696 78752 144702 78804
rect 146110 78752 146116 78804
rect 146168 78792 146174 78804
rect 148502 78792 148508 78804
rect 146168 78764 148508 78792
rect 146168 78752 146174 78764
rect 148502 78752 148508 78764
rect 148560 78752 148566 78804
rect 172330 78752 172336 78804
rect 172388 78792 172394 78804
rect 217134 78792 217140 78804
rect 172388 78764 217140 78792
rect 172388 78752 172394 78764
rect 217134 78752 217140 78764
rect 217192 78752 217198 78804
rect 129642 78684 129648 78736
rect 129700 78724 129706 78736
rect 138014 78724 138020 78736
rect 129700 78696 138020 78724
rect 129700 78684 129706 78696
rect 138014 78684 138020 78696
rect 138072 78684 138078 78736
rect 168374 78684 168380 78736
rect 168432 78724 168438 78736
rect 172054 78724 172060 78736
rect 168432 78696 172060 78724
rect 168432 78684 168438 78696
rect 172054 78684 172060 78696
rect 172112 78684 172118 78736
rect 181346 78684 181352 78736
rect 181404 78724 181410 78736
rect 182174 78724 182180 78736
rect 181404 78696 182180 78724
rect 181404 78684 181410 78696
rect 182174 78684 182180 78696
rect 182232 78684 182238 78736
rect 120994 78616 121000 78668
rect 121052 78656 121058 78668
rect 135806 78656 135812 78668
rect 121052 78628 135812 78656
rect 121052 78616 121058 78628
rect 135806 78616 135812 78628
rect 135864 78616 135870 78668
rect 136634 78616 136640 78668
rect 136692 78656 136698 78668
rect 143258 78656 143264 78668
rect 136692 78628 143264 78656
rect 136692 78616 136698 78628
rect 143258 78616 143264 78628
rect 143316 78616 143322 78668
rect 154574 78616 154580 78668
rect 154632 78656 154638 78668
rect 154942 78656 154948 78668
rect 154632 78628 154948 78656
rect 154632 78616 154638 78628
rect 154942 78616 154948 78628
rect 155000 78616 155006 78668
rect 155586 78616 155592 78668
rect 155644 78656 155650 78668
rect 158346 78656 158352 78668
rect 155644 78628 158352 78656
rect 155644 78616 155650 78628
rect 158346 78616 158352 78628
rect 158404 78616 158410 78668
rect 160094 78616 160100 78668
rect 160152 78656 160158 78668
rect 160278 78656 160284 78668
rect 160152 78628 160284 78656
rect 160152 78616 160158 78628
rect 160278 78616 160284 78628
rect 160336 78616 160342 78668
rect 168650 78616 168656 78668
rect 168708 78656 168714 78668
rect 169294 78656 169300 78668
rect 168708 78628 169300 78656
rect 168708 78616 168714 78628
rect 169294 78616 169300 78628
rect 169352 78616 169358 78668
rect 174078 78616 174084 78668
rect 174136 78656 174142 78668
rect 188798 78656 188804 78668
rect 174136 78628 188804 78656
rect 174136 78616 174142 78628
rect 188798 78616 188804 78628
rect 188856 78616 188862 78668
rect 131022 78548 131028 78600
rect 131080 78588 131086 78600
rect 138382 78588 138388 78600
rect 131080 78560 138388 78588
rect 131080 78548 131086 78560
rect 138382 78548 138388 78560
rect 138440 78548 138446 78600
rect 142614 78548 142620 78600
rect 142672 78588 142678 78600
rect 142798 78588 142804 78600
rect 142672 78560 142804 78588
rect 142672 78548 142678 78560
rect 142798 78548 142804 78560
rect 142856 78548 142862 78600
rect 166994 78548 167000 78600
rect 167052 78588 167058 78600
rect 168190 78588 168196 78600
rect 167052 78560 168196 78588
rect 167052 78548 167058 78560
rect 168190 78548 168196 78560
rect 168248 78548 168254 78600
rect 173066 78548 173072 78600
rect 173124 78588 173130 78600
rect 209958 78588 209964 78600
rect 173124 78560 209964 78588
rect 173124 78548 173130 78560
rect 209958 78548 209964 78560
rect 210016 78548 210022 78600
rect 104526 78480 104532 78532
rect 104584 78520 104590 78532
rect 127434 78520 127440 78532
rect 104584 78492 127440 78520
rect 104584 78480 104590 78492
rect 127434 78480 127440 78492
rect 127492 78480 127498 78532
rect 131850 78480 131856 78532
rect 131908 78520 131914 78532
rect 141510 78520 141516 78532
rect 131908 78492 141516 78520
rect 131908 78480 131914 78492
rect 141510 78480 141516 78492
rect 141568 78480 141574 78532
rect 175918 78480 175924 78532
rect 175976 78520 175982 78532
rect 207842 78520 207848 78532
rect 175976 78492 207848 78520
rect 175976 78480 175982 78492
rect 207842 78480 207848 78492
rect 207900 78480 207906 78532
rect 104066 78412 104072 78464
rect 104124 78452 104130 78464
rect 129642 78452 129648 78464
rect 104124 78424 129648 78452
rect 104124 78412 104130 78424
rect 129642 78412 129648 78424
rect 129700 78412 129706 78464
rect 131114 78412 131120 78464
rect 131172 78452 131178 78464
rect 132310 78452 132316 78464
rect 131172 78424 132316 78452
rect 131172 78412 131178 78424
rect 132310 78412 132316 78424
rect 132368 78412 132374 78464
rect 132494 78412 132500 78464
rect 132552 78452 132558 78464
rect 136726 78452 136732 78464
rect 132552 78424 136732 78452
rect 132552 78412 132558 78424
rect 136726 78412 136732 78424
rect 136784 78412 136790 78464
rect 155862 78412 155868 78464
rect 155920 78452 155926 78464
rect 156598 78452 156604 78464
rect 155920 78424 156604 78452
rect 155920 78412 155926 78424
rect 156598 78412 156604 78424
rect 156656 78412 156662 78464
rect 166534 78412 166540 78464
rect 166592 78452 166598 78464
rect 166592 78424 168374 78452
rect 166592 78412 166598 78424
rect 104434 78344 104440 78396
rect 104492 78384 104498 78396
rect 128538 78384 128544 78396
rect 104492 78356 128544 78384
rect 104492 78344 104498 78356
rect 128538 78344 128544 78356
rect 128596 78344 128602 78396
rect 131206 78344 131212 78396
rect 131264 78384 131270 78396
rect 138934 78384 138940 78396
rect 131264 78356 138940 78384
rect 131264 78344 131270 78356
rect 138934 78344 138940 78356
rect 138992 78344 138998 78396
rect 140406 78344 140412 78396
rect 140464 78384 140470 78396
rect 147398 78384 147404 78396
rect 140464 78356 147404 78384
rect 140464 78344 140470 78356
rect 147398 78344 147404 78356
rect 147456 78344 147462 78396
rect 163222 78344 163228 78396
rect 163280 78384 163286 78396
rect 166626 78384 166632 78396
rect 163280 78356 166632 78384
rect 163280 78344 163286 78356
rect 166626 78344 166632 78356
rect 166684 78344 166690 78396
rect 168346 78384 168374 78424
rect 171778 78412 171784 78464
rect 171836 78452 171842 78464
rect 206186 78452 206192 78464
rect 171836 78424 206192 78452
rect 171836 78412 171842 78424
rect 206186 78412 206192 78424
rect 206244 78412 206250 78464
rect 188890 78384 188896 78396
rect 168346 78356 188896 78384
rect 188890 78344 188896 78356
rect 188948 78344 188954 78396
rect 106826 78276 106832 78328
rect 106884 78316 106890 78328
rect 131298 78316 131304 78328
rect 106884 78288 131304 78316
rect 106884 78276 106890 78288
rect 131298 78276 131304 78288
rect 131356 78276 131362 78328
rect 149974 78316 149980 78328
rect 137986 78288 149980 78316
rect 122282 78208 122288 78260
rect 122340 78248 122346 78260
rect 135438 78248 135444 78260
rect 122340 78220 135444 78248
rect 122340 78208 122346 78220
rect 135438 78208 135444 78220
rect 135496 78208 135502 78260
rect 121270 78140 121276 78192
rect 121328 78180 121334 78192
rect 133690 78180 133696 78192
rect 121328 78152 133696 78180
rect 121328 78140 121334 78152
rect 133690 78140 133696 78152
rect 133748 78140 133754 78192
rect 106918 78072 106924 78124
rect 106976 78112 106982 78124
rect 125226 78112 125232 78124
rect 106976 78084 125232 78112
rect 106976 78072 106982 78084
rect 125226 78072 125232 78084
rect 125284 78072 125290 78124
rect 132310 78072 132316 78124
rect 132368 78112 132374 78124
rect 137986 78112 138014 78288
rect 149974 78276 149980 78288
rect 150032 78276 150038 78328
rect 152458 78276 152464 78328
rect 152516 78316 152522 78328
rect 162302 78316 162308 78328
rect 152516 78288 162308 78316
rect 152516 78276 152522 78288
rect 162302 78276 162308 78288
rect 162360 78276 162366 78328
rect 163130 78276 163136 78328
rect 163188 78316 163194 78328
rect 165522 78316 165528 78328
rect 163188 78288 165528 78316
rect 163188 78276 163194 78288
rect 165522 78276 165528 78288
rect 165580 78276 165586 78328
rect 168558 78276 168564 78328
rect 168616 78316 168622 78328
rect 169386 78316 169392 78328
rect 168616 78288 169392 78316
rect 168616 78276 168622 78288
rect 169386 78276 169392 78288
rect 169444 78276 169450 78328
rect 169662 78276 169668 78328
rect 169720 78316 169726 78328
rect 188706 78316 188712 78328
rect 169720 78288 188712 78316
rect 169720 78276 169726 78288
rect 188706 78276 188712 78288
rect 188764 78276 188770 78328
rect 138934 78208 138940 78260
rect 138992 78248 138998 78260
rect 142246 78248 142252 78260
rect 138992 78220 142252 78248
rect 138992 78208 138998 78220
rect 142246 78208 142252 78220
rect 142304 78208 142310 78260
rect 148870 78208 148876 78260
rect 148928 78248 148934 78260
rect 158162 78248 158168 78260
rect 148928 78220 158168 78248
rect 148928 78208 148934 78220
rect 158162 78208 158168 78220
rect 158220 78208 158226 78260
rect 161198 78208 161204 78260
rect 161256 78248 161262 78260
rect 161256 78220 166120 78248
rect 161256 78208 161262 78220
rect 157242 78140 157248 78192
rect 157300 78180 157306 78192
rect 165982 78180 165988 78192
rect 157300 78152 165988 78180
rect 157300 78140 157306 78152
rect 165982 78140 165988 78152
rect 166040 78140 166046 78192
rect 166092 78180 166120 78220
rect 167270 78208 167276 78260
rect 167328 78248 167334 78260
rect 177390 78248 177396 78260
rect 167328 78220 177396 78248
rect 167328 78208 167334 78220
rect 177390 78208 177396 78220
rect 177448 78208 177454 78260
rect 181806 78208 181812 78260
rect 181864 78248 181870 78260
rect 181864 78220 190454 78248
rect 181864 78208 181870 78220
rect 169478 78180 169484 78192
rect 166092 78152 169484 78180
rect 169478 78140 169484 78152
rect 169536 78140 169542 78192
rect 172974 78140 172980 78192
rect 173032 78180 173038 78192
rect 174722 78180 174728 78192
rect 173032 78152 174728 78180
rect 173032 78140 173038 78152
rect 174722 78140 174728 78152
rect 174780 78140 174786 78192
rect 174814 78140 174820 78192
rect 174872 78180 174878 78192
rect 174998 78180 175004 78192
rect 174872 78152 175004 78180
rect 174872 78140 174878 78152
rect 174998 78140 175004 78152
rect 175056 78180 175062 78192
rect 189718 78180 189724 78192
rect 175056 78152 189724 78180
rect 175056 78140 175062 78152
rect 189718 78140 189724 78152
rect 189776 78140 189782 78192
rect 190426 78180 190454 78220
rect 195238 78180 195244 78192
rect 190426 78152 195244 78180
rect 195238 78140 195244 78152
rect 195296 78140 195302 78192
rect 148778 78112 148784 78124
rect 132368 78084 138014 78112
rect 142816 78084 148784 78112
rect 132368 78072 132374 78084
rect 107470 78004 107476 78056
rect 107528 78044 107534 78056
rect 128446 78044 128452 78056
rect 107528 78016 128452 78044
rect 107528 78004 107534 78016
rect 128446 78004 128452 78016
rect 128504 78004 128510 78056
rect 128998 78004 129004 78056
rect 129056 78044 129062 78056
rect 134242 78044 134248 78056
rect 129056 78016 134248 78044
rect 129056 78004 129062 78016
rect 134242 78004 134248 78016
rect 134300 78004 134306 78056
rect 136726 78004 136732 78056
rect 136784 78044 136790 78056
rect 142816 78044 142844 78084
rect 148778 78072 148784 78084
rect 148836 78072 148842 78124
rect 153378 78072 153384 78124
rect 153436 78112 153442 78124
rect 154114 78112 154120 78124
rect 153436 78084 154120 78112
rect 153436 78072 153442 78084
rect 154114 78072 154120 78084
rect 154172 78072 154178 78124
rect 158162 78072 158168 78124
rect 158220 78112 158226 78124
rect 158806 78112 158812 78124
rect 158220 78084 158812 78112
rect 158220 78072 158226 78084
rect 158806 78072 158812 78084
rect 158864 78072 158870 78124
rect 160370 78072 160376 78124
rect 160428 78112 160434 78124
rect 166166 78112 166172 78124
rect 160428 78084 166172 78112
rect 160428 78072 160434 78084
rect 166166 78072 166172 78084
rect 166224 78072 166230 78124
rect 167454 78072 167460 78124
rect 167512 78112 167518 78124
rect 182082 78112 182088 78124
rect 167512 78084 182088 78112
rect 167512 78072 167518 78084
rect 182082 78072 182088 78084
rect 182140 78072 182146 78124
rect 182910 78072 182916 78124
rect 182968 78112 182974 78124
rect 196802 78112 196808 78124
rect 182968 78084 196808 78112
rect 182968 78072 182974 78084
rect 196802 78072 196808 78084
rect 196860 78072 196866 78124
rect 155678 78044 155684 78056
rect 136784 78016 142844 78044
rect 147646 78016 155684 78044
rect 136784 78004 136790 78016
rect 103974 77936 103980 77988
rect 104032 77976 104038 77988
rect 104032 77948 128354 77976
rect 104032 77936 104038 77948
rect 128326 77840 128354 77948
rect 135898 77936 135904 77988
rect 135956 77976 135962 77988
rect 147646 77976 147674 78016
rect 155678 78004 155684 78016
rect 155736 78004 155742 78056
rect 157886 78004 157892 78056
rect 157944 78044 157950 78056
rect 169662 78044 169668 78056
rect 157944 78016 169668 78044
rect 157944 78004 157950 78016
rect 169662 78004 169668 78016
rect 169720 78004 169726 78056
rect 170490 78004 170496 78056
rect 170548 78044 170554 78056
rect 180518 78044 180524 78056
rect 170548 78016 180524 78044
rect 170548 78004 170554 78016
rect 180518 78004 180524 78016
rect 180576 78004 180582 78056
rect 180702 78004 180708 78056
rect 180760 78044 180766 78056
rect 204990 78044 204996 78056
rect 180760 78016 204996 78044
rect 180760 78004 180766 78016
rect 204990 78004 204996 78016
rect 205048 78004 205054 78056
rect 135956 77948 147674 77976
rect 135956 77936 135962 77948
rect 148318 77936 148324 77988
rect 148376 77976 148382 77988
rect 148962 77976 148968 77988
rect 148376 77948 148968 77976
rect 148376 77936 148382 77948
rect 148962 77936 148968 77948
rect 149020 77936 149026 77988
rect 156506 77936 156512 77988
rect 156564 77976 156570 77988
rect 169294 77976 169300 77988
rect 156564 77948 169300 77976
rect 156564 77936 156570 77948
rect 169294 77936 169300 77948
rect 169352 77936 169358 77988
rect 180334 77936 180340 77988
rect 180392 77976 180398 77988
rect 206370 77976 206376 77988
rect 180392 77948 206376 77976
rect 180392 77936 180398 77948
rect 206370 77936 206376 77948
rect 206428 77936 206434 77988
rect 137370 77868 137376 77920
rect 137428 77908 137434 77920
rect 140498 77908 140504 77920
rect 137428 77880 140504 77908
rect 137428 77868 137434 77880
rect 140498 77868 140504 77880
rect 140556 77868 140562 77920
rect 154022 77908 154028 77920
rect 144886 77880 154028 77908
rect 137922 77840 137928 77852
rect 128326 77812 137928 77840
rect 137922 77800 137928 77812
rect 137980 77800 137986 77852
rect 138382 77800 138388 77852
rect 138440 77840 138446 77852
rect 138566 77840 138572 77852
rect 138440 77812 138572 77840
rect 138440 77800 138446 77812
rect 138566 77800 138572 77812
rect 138624 77800 138630 77852
rect 141418 77800 141424 77852
rect 141476 77840 141482 77852
rect 144362 77840 144368 77852
rect 141476 77812 144368 77840
rect 141476 77800 141482 77812
rect 144362 77800 144368 77812
rect 144420 77800 144426 77852
rect 96246 77732 96252 77784
rect 96304 77772 96310 77784
rect 138842 77772 138848 77784
rect 96304 77744 138848 77772
rect 96304 77732 96310 77744
rect 138842 77732 138848 77744
rect 138900 77732 138906 77784
rect 122006 77664 122012 77716
rect 122064 77704 122070 77716
rect 135070 77704 135076 77716
rect 122064 77676 135076 77704
rect 122064 77664 122070 77676
rect 135070 77664 135076 77676
rect 135128 77704 135134 77716
rect 144886 77704 144914 77880
rect 154022 77868 154028 77880
rect 154080 77868 154086 77920
rect 163222 77868 163228 77920
rect 163280 77908 163286 77920
rect 163958 77908 163964 77920
rect 163280 77880 163964 77908
rect 163280 77868 163286 77880
rect 163958 77868 163964 77880
rect 164016 77868 164022 77920
rect 167270 77868 167276 77920
rect 167328 77908 167334 77920
rect 167546 77908 167552 77920
rect 167328 77880 167552 77908
rect 167328 77868 167334 77880
rect 167546 77868 167552 77880
rect 167604 77868 167610 77920
rect 170950 77868 170956 77920
rect 171008 77908 171014 77920
rect 173526 77908 173532 77920
rect 171008 77880 173532 77908
rect 171008 77868 171014 77880
rect 173526 77868 173532 77880
rect 173584 77868 173590 77920
rect 182818 77868 182824 77920
rect 182876 77908 182882 77920
rect 195606 77908 195612 77920
rect 182876 77880 195612 77908
rect 182876 77868 182882 77880
rect 195606 77868 195612 77880
rect 195664 77868 195670 77920
rect 147766 77800 147772 77852
rect 147824 77840 147830 77852
rect 148594 77840 148600 77852
rect 147824 77812 148600 77840
rect 147824 77800 147830 77812
rect 148594 77800 148600 77812
rect 148652 77800 148658 77852
rect 157702 77732 157708 77784
rect 157760 77772 157766 77784
rect 212994 77772 213000 77784
rect 157760 77744 213000 77772
rect 157760 77732 157766 77744
rect 212994 77732 213000 77744
rect 213052 77732 213058 77784
rect 135128 77676 144914 77704
rect 135128 77664 135134 77676
rect 165798 77664 165804 77716
rect 165856 77704 165862 77716
rect 166350 77704 166356 77716
rect 165856 77676 166356 77704
rect 165856 77664 165862 77676
rect 166350 77664 166356 77676
rect 166408 77664 166414 77716
rect 167914 77664 167920 77716
rect 167972 77704 167978 77716
rect 169018 77704 169024 77716
rect 167972 77676 169024 77704
rect 167972 77664 167978 77676
rect 169018 77664 169024 77676
rect 169076 77664 169082 77716
rect 170306 77664 170312 77716
rect 170364 77704 170370 77716
rect 189902 77704 189908 77716
rect 170364 77676 189908 77704
rect 170364 77664 170370 77676
rect 189902 77664 189908 77676
rect 189960 77664 189966 77716
rect 122806 77608 131114 77636
rect 99098 77528 99104 77580
rect 99156 77568 99162 77580
rect 122806 77568 122834 77608
rect 99156 77540 122834 77568
rect 131086 77568 131114 77608
rect 138566 77596 138572 77648
rect 138624 77636 138630 77648
rect 140314 77636 140320 77648
rect 138624 77608 140320 77636
rect 138624 77596 138630 77608
rect 140314 77596 140320 77608
rect 140372 77636 140378 77648
rect 140372 77608 147674 77636
rect 140372 77596 140378 77608
rect 139946 77568 139952 77580
rect 131086 77540 139952 77568
rect 99156 77528 99162 77540
rect 139946 77528 139952 77540
rect 140004 77528 140010 77580
rect 140590 77528 140596 77580
rect 140648 77568 140654 77580
rect 144822 77568 144828 77580
rect 140648 77540 144828 77568
rect 140648 77528 140654 77540
rect 144822 77528 144828 77540
rect 144880 77528 144886 77580
rect 138750 77460 138756 77512
rect 138808 77500 138814 77512
rect 146294 77500 146300 77512
rect 138808 77472 146300 77500
rect 138808 77460 138814 77472
rect 146294 77460 146300 77472
rect 146352 77460 146358 77512
rect 134150 77324 134156 77376
rect 134208 77364 134214 77376
rect 134886 77364 134892 77376
rect 134208 77336 134892 77364
rect 134208 77324 134214 77336
rect 134886 77324 134892 77336
rect 134944 77324 134950 77376
rect 132126 77256 132132 77308
rect 132184 77296 132190 77308
rect 139118 77296 139124 77308
rect 132184 77268 139124 77296
rect 132184 77256 132190 77268
rect 139118 77256 139124 77268
rect 139176 77256 139182 77308
rect 147646 77296 147674 77608
rect 163590 77596 163596 77648
rect 163648 77636 163654 77648
rect 170950 77636 170956 77648
rect 163648 77608 170956 77636
rect 163648 77596 163654 77608
rect 170950 77596 170956 77608
rect 171008 77596 171014 77648
rect 147766 77528 147772 77580
rect 147824 77568 147830 77580
rect 148686 77568 148692 77580
rect 147824 77540 148692 77568
rect 147824 77528 147830 77540
rect 148686 77528 148692 77540
rect 148744 77528 148750 77580
rect 165062 77460 165068 77512
rect 165120 77500 165126 77512
rect 172514 77500 172520 77512
rect 165120 77472 172520 77500
rect 165120 77460 165126 77472
rect 172514 77460 172520 77472
rect 172572 77460 172578 77512
rect 156874 77296 156880 77308
rect 147646 77268 156880 77296
rect 156874 77256 156880 77268
rect 156932 77256 156938 77308
rect 159450 77256 159456 77308
rect 159508 77296 159514 77308
rect 163866 77296 163872 77308
rect 159508 77268 163872 77296
rect 159508 77256 159514 77268
rect 163866 77256 163872 77268
rect 163924 77256 163930 77308
rect 2774 77188 2780 77240
rect 2832 77228 2838 77240
rect 4798 77228 4804 77240
rect 2832 77200 4804 77228
rect 2832 77188 2838 77200
rect 4798 77188 4804 77200
rect 4856 77188 4862 77240
rect 120074 77188 120080 77240
rect 120132 77228 120138 77240
rect 142338 77228 142344 77240
rect 120132 77200 142344 77228
rect 120132 77188 120138 77200
rect 142338 77188 142344 77200
rect 142396 77188 142402 77240
rect 158622 77188 158628 77240
rect 158680 77228 158686 77240
rect 160554 77228 160560 77240
rect 158680 77200 160560 77228
rect 158680 77188 158686 77200
rect 160554 77188 160560 77200
rect 160612 77188 160618 77240
rect 176102 77188 176108 77240
rect 176160 77228 176166 77240
rect 200482 77228 200488 77240
rect 176160 77200 200488 77228
rect 176160 77188 176166 77200
rect 200482 77188 200488 77200
rect 200540 77188 200546 77240
rect 115290 77120 115296 77172
rect 115348 77160 115354 77172
rect 115348 77132 128354 77160
rect 115348 77120 115354 77132
rect 128326 77092 128354 77132
rect 140038 77120 140044 77172
rect 140096 77160 140102 77172
rect 140222 77160 140228 77172
rect 140096 77132 140228 77160
rect 140096 77120 140102 77132
rect 140222 77120 140228 77132
rect 140280 77120 140286 77172
rect 152918 77120 152924 77172
rect 152976 77160 152982 77172
rect 215570 77160 215576 77172
rect 152976 77132 215576 77160
rect 152976 77120 152982 77132
rect 215570 77120 215576 77132
rect 215628 77120 215634 77172
rect 140406 77092 140412 77104
rect 128326 77064 140412 77092
rect 140406 77052 140412 77064
rect 140464 77052 140470 77104
rect 141694 77052 141700 77104
rect 141752 77092 141758 77104
rect 143074 77092 143080 77104
rect 141752 77064 143080 77092
rect 141752 77052 141758 77064
rect 143074 77052 143080 77064
rect 143132 77052 143138 77104
rect 159266 77052 159272 77104
rect 159324 77092 159330 77104
rect 159450 77092 159456 77104
rect 159324 77064 159456 77092
rect 159324 77052 159330 77064
rect 159450 77052 159456 77064
rect 159508 77052 159514 77104
rect 172422 77052 172428 77104
rect 172480 77092 172486 77104
rect 211890 77092 211896 77104
rect 172480 77064 211896 77092
rect 172480 77052 172486 77064
rect 211890 77052 211896 77064
rect 211948 77052 211954 77104
rect 117774 76984 117780 77036
rect 117832 77024 117838 77036
rect 166534 77024 166540 77036
rect 117832 76996 166540 77024
rect 117832 76984 117838 76996
rect 166534 76984 166540 76996
rect 166592 76984 166598 77036
rect 173618 76984 173624 77036
rect 173676 77024 173682 77036
rect 211798 77024 211804 77036
rect 173676 76996 211804 77024
rect 173676 76984 173682 76996
rect 211798 76984 211804 76996
rect 211856 76984 211862 77036
rect 115842 76916 115848 76968
rect 115900 76956 115906 76968
rect 142614 76956 142620 76968
rect 115900 76928 142620 76956
rect 115900 76916 115906 76928
rect 142614 76916 142620 76928
rect 142672 76916 142678 76968
rect 156046 76916 156052 76968
rect 156104 76956 156110 76968
rect 157702 76956 157708 76968
rect 156104 76928 157708 76956
rect 156104 76916 156110 76928
rect 157702 76916 157708 76928
rect 157760 76916 157766 76968
rect 175366 76916 175372 76968
rect 175424 76956 175430 76968
rect 218422 76956 218428 76968
rect 175424 76928 218428 76956
rect 175424 76916 175430 76928
rect 218422 76916 218428 76928
rect 218480 76916 218486 76968
rect 114094 76848 114100 76900
rect 114152 76888 114158 76900
rect 146110 76888 146116 76900
rect 114152 76860 146116 76888
rect 114152 76848 114158 76860
rect 146110 76848 146116 76860
rect 146168 76848 146174 76900
rect 156414 76848 156420 76900
rect 156472 76888 156478 76900
rect 158714 76888 158720 76900
rect 156472 76860 158720 76888
rect 156472 76848 156478 76860
rect 158714 76848 158720 76860
rect 158772 76888 158778 76900
rect 192478 76888 192484 76900
rect 158772 76860 192484 76888
rect 158772 76848 158778 76860
rect 192478 76848 192484 76860
rect 192536 76848 192542 76900
rect 113726 76780 113732 76832
rect 113784 76820 113790 76832
rect 147582 76820 147588 76832
rect 113784 76792 147588 76820
rect 113784 76780 113790 76792
rect 147582 76780 147588 76792
rect 147640 76780 147646 76832
rect 172790 76780 172796 76832
rect 172848 76820 172854 76832
rect 208946 76820 208952 76832
rect 172848 76792 208952 76820
rect 172848 76780 172854 76792
rect 208946 76780 208952 76792
rect 209004 76780 209010 76832
rect 118326 76712 118332 76764
rect 118384 76752 118390 76764
rect 149238 76752 149244 76764
rect 118384 76724 149244 76752
rect 118384 76712 118390 76724
rect 149238 76712 149244 76724
rect 149296 76752 149302 76764
rect 149296 76724 157334 76752
rect 149296 76712 149302 76724
rect 119338 76644 119344 76696
rect 119396 76684 119402 76696
rect 149606 76684 149612 76696
rect 119396 76656 149612 76684
rect 119396 76644 119402 76656
rect 149606 76644 149612 76656
rect 149664 76644 149670 76696
rect 94958 76576 94964 76628
rect 95016 76616 95022 76628
rect 129642 76616 129648 76628
rect 95016 76588 129648 76616
rect 95016 76576 95022 76588
rect 129642 76576 129648 76588
rect 129700 76576 129706 76628
rect 135622 76576 135628 76628
rect 135680 76616 135686 76628
rect 136082 76616 136088 76628
rect 135680 76588 136088 76616
rect 135680 76576 135686 76588
rect 136082 76576 136088 76588
rect 136140 76576 136146 76628
rect 139578 76576 139584 76628
rect 139636 76616 139642 76628
rect 139854 76616 139860 76628
rect 139636 76588 139860 76616
rect 139636 76576 139642 76588
rect 139854 76576 139860 76588
rect 139912 76576 139918 76628
rect 141326 76576 141332 76628
rect 141384 76616 141390 76628
rect 141694 76616 141700 76628
rect 141384 76588 141700 76616
rect 141384 76576 141390 76588
rect 141694 76576 141700 76588
rect 141752 76576 141758 76628
rect 142614 76576 142620 76628
rect 142672 76616 142678 76628
rect 145006 76616 145012 76628
rect 142672 76588 145012 76616
rect 142672 76576 142678 76588
rect 145006 76576 145012 76588
rect 145064 76576 145070 76628
rect 153746 76576 153752 76628
rect 153804 76616 153810 76628
rect 154482 76616 154488 76628
rect 153804 76588 154488 76616
rect 153804 76576 153810 76588
rect 154482 76576 154488 76588
rect 154540 76576 154546 76628
rect 154666 76576 154672 76628
rect 154724 76616 154730 76628
rect 154850 76616 154856 76628
rect 154724 76588 154856 76616
rect 154724 76576 154730 76588
rect 154850 76576 154856 76588
rect 154908 76576 154914 76628
rect 156506 76576 156512 76628
rect 156564 76616 156570 76628
rect 156966 76616 156972 76628
rect 156564 76588 156972 76616
rect 156564 76576 156570 76588
rect 156966 76576 156972 76588
rect 157024 76576 157030 76628
rect 67634 76508 67640 76560
rect 67692 76548 67698 76560
rect 115198 76548 115204 76560
rect 67692 76520 115204 76548
rect 67692 76508 67698 76520
rect 115198 76508 115204 76520
rect 115256 76548 115262 76560
rect 115842 76548 115848 76560
rect 115256 76520 115848 76548
rect 115256 76508 115262 76520
rect 115842 76508 115848 76520
rect 115900 76508 115906 76560
rect 135530 76508 135536 76560
rect 135588 76548 135594 76560
rect 136358 76548 136364 76560
rect 135588 76520 136364 76548
rect 135588 76508 135594 76520
rect 136358 76508 136364 76520
rect 136416 76508 136422 76560
rect 157306 76548 157334 76724
rect 177482 76712 177488 76764
rect 177540 76752 177546 76764
rect 209958 76752 209964 76764
rect 177540 76724 209964 76752
rect 177540 76712 177546 76724
rect 209958 76712 209964 76724
rect 210016 76712 210022 76764
rect 168466 76644 168472 76696
rect 168524 76684 168530 76696
rect 203334 76684 203340 76696
rect 168524 76656 203340 76684
rect 168524 76644 168530 76656
rect 203334 76644 203340 76656
rect 203392 76644 203398 76696
rect 165706 76576 165712 76628
rect 165764 76616 165770 76628
rect 176470 76616 176476 76628
rect 165764 76588 176476 76616
rect 165764 76576 165770 76588
rect 176470 76576 176476 76588
rect 176528 76576 176534 76628
rect 179782 76576 179788 76628
rect 179840 76616 179846 76628
rect 203058 76616 203064 76628
rect 179840 76588 203064 76616
rect 179840 76576 179846 76588
rect 203058 76576 203064 76588
rect 203116 76576 203122 76628
rect 289814 76548 289820 76560
rect 157306 76520 289820 76548
rect 289814 76508 289820 76520
rect 289872 76508 289878 76560
rect 102134 76440 102140 76492
rect 102192 76480 102198 76492
rect 133138 76480 133144 76492
rect 102192 76452 133144 76480
rect 102192 76440 102198 76452
rect 133138 76440 133144 76452
rect 133196 76440 133202 76492
rect 141050 76440 141056 76492
rect 141108 76480 141114 76492
rect 141786 76480 141792 76492
rect 141108 76452 141792 76480
rect 141108 76440 141114 76452
rect 141786 76440 141792 76452
rect 141844 76440 141850 76492
rect 155310 76440 155316 76492
rect 155368 76480 155374 76492
rect 158530 76480 158536 76492
rect 155368 76452 158536 76480
rect 155368 76440 155374 76452
rect 158530 76440 158536 76452
rect 158588 76440 158594 76492
rect 165706 76440 165712 76492
rect 165764 76480 165770 76492
rect 166810 76480 166816 76492
rect 165764 76452 166816 76480
rect 165764 76440 165770 76452
rect 166810 76440 166816 76452
rect 166868 76440 166874 76492
rect 119154 76372 119160 76424
rect 119212 76412 119218 76424
rect 156414 76412 156420 76424
rect 119212 76384 156420 76412
rect 119212 76372 119218 76384
rect 156414 76372 156420 76384
rect 156472 76372 156478 76424
rect 165522 76372 165528 76424
rect 165580 76412 165586 76424
rect 204806 76412 204812 76424
rect 165580 76384 204812 76412
rect 165580 76372 165586 76384
rect 204806 76372 204812 76384
rect 204864 76372 204870 76424
rect 94682 76304 94688 76356
rect 94740 76344 94746 76356
rect 163498 76344 163504 76356
rect 94740 76316 163504 76344
rect 94740 76304 94746 76316
rect 163498 76304 163504 76316
rect 163556 76304 163562 76356
rect 180334 76344 180340 76356
rect 166736 76316 180340 76344
rect 113634 76236 113640 76288
rect 113692 76276 113698 76288
rect 166442 76276 166448 76288
rect 113692 76248 166448 76276
rect 113692 76236 113698 76248
rect 166442 76236 166448 76248
rect 166500 76276 166506 76288
rect 166736 76276 166764 76316
rect 180334 76304 180340 76316
rect 180392 76304 180398 76356
rect 166500 76248 166764 76276
rect 166500 76236 166506 76248
rect 170030 76236 170036 76288
rect 170088 76276 170094 76288
rect 180702 76276 180708 76288
rect 170088 76248 180708 76276
rect 170088 76236 170094 76248
rect 180702 76236 180708 76248
rect 180760 76236 180766 76288
rect 135714 76168 135720 76220
rect 135772 76208 135778 76220
rect 136450 76208 136456 76220
rect 135772 76180 136456 76208
rect 135772 76168 135778 76180
rect 136450 76168 136456 76180
rect 136508 76168 136514 76220
rect 140958 76168 140964 76220
rect 141016 76208 141022 76220
rect 141602 76208 141608 76220
rect 141016 76180 141608 76208
rect 141016 76168 141022 76180
rect 141602 76168 141608 76180
rect 141660 76168 141666 76220
rect 155126 76168 155132 76220
rect 155184 76208 155190 76220
rect 155586 76208 155592 76220
rect 155184 76180 155592 76208
rect 155184 76168 155190 76180
rect 155586 76168 155592 76180
rect 155644 76168 155650 76220
rect 156414 76168 156420 76220
rect 156472 76208 156478 76220
rect 156598 76208 156604 76220
rect 156472 76180 156604 76208
rect 156472 76168 156478 76180
rect 156598 76168 156604 76180
rect 156656 76168 156662 76220
rect 158254 76168 158260 76220
rect 158312 76208 158318 76220
rect 158714 76208 158720 76220
rect 158312 76180 158720 76208
rect 158312 76168 158318 76180
rect 158714 76168 158720 76180
rect 158772 76168 158778 76220
rect 159082 76168 159088 76220
rect 159140 76208 159146 76220
rect 159358 76208 159364 76220
rect 159140 76180 159364 76208
rect 159140 76168 159146 76180
rect 159358 76168 159364 76180
rect 159416 76168 159422 76220
rect 166258 76168 166264 76220
rect 166316 76208 166322 76220
rect 166902 76208 166908 76220
rect 166316 76180 166908 76208
rect 166316 76168 166322 76180
rect 166902 76168 166908 76180
rect 166960 76168 166966 76220
rect 132678 76100 132684 76152
rect 132736 76140 132742 76152
rect 132862 76140 132868 76152
rect 132736 76112 132868 76140
rect 132736 76100 132742 76112
rect 132862 76100 132868 76112
rect 132920 76100 132926 76152
rect 136174 76100 136180 76152
rect 136232 76140 136238 76152
rect 136542 76140 136548 76152
rect 136232 76112 136548 76140
rect 136232 76100 136238 76112
rect 136542 76100 136548 76112
rect 136600 76100 136606 76152
rect 154942 76100 154948 76152
rect 155000 76140 155006 76152
rect 155402 76140 155408 76152
rect 155000 76112 155408 76140
rect 155000 76100 155006 76112
rect 155402 76100 155408 76112
rect 155460 76100 155466 76152
rect 156230 76100 156236 76152
rect 156288 76140 156294 76152
rect 157334 76140 157340 76152
rect 156288 76112 157340 76140
rect 156288 76100 156294 76112
rect 157334 76100 157340 76112
rect 157392 76100 157398 76152
rect 175182 76100 175188 76152
rect 175240 76140 175246 76152
rect 177942 76140 177948 76152
rect 175240 76112 177948 76140
rect 175240 76100 175246 76112
rect 177942 76100 177948 76112
rect 178000 76100 178006 76152
rect 135346 76032 135352 76084
rect 135404 76072 135410 76084
rect 136450 76072 136456 76084
rect 135404 76044 136456 76072
rect 135404 76032 135410 76044
rect 136450 76032 136456 76044
rect 136508 76032 136514 76084
rect 136818 76032 136824 76084
rect 136876 76072 136882 76084
rect 137278 76072 137284 76084
rect 136876 76044 137284 76072
rect 136876 76032 136882 76044
rect 137278 76032 137284 76044
rect 137336 76032 137342 76084
rect 138014 76032 138020 76084
rect 138072 76072 138078 76084
rect 139026 76072 139032 76084
rect 138072 76044 139032 76072
rect 138072 76032 138078 76044
rect 139026 76032 139032 76044
rect 139084 76032 139090 76084
rect 158990 76032 158996 76084
rect 159048 76072 159054 76084
rect 159358 76072 159364 76084
rect 159048 76044 159364 76072
rect 159048 76032 159054 76044
rect 159358 76032 159364 76044
rect 159416 76032 159422 76084
rect 161750 76032 161756 76084
rect 161808 76072 161814 76084
rect 166258 76072 166264 76084
rect 161808 76044 166264 76072
rect 161808 76032 161814 76044
rect 166258 76032 166264 76044
rect 166316 76032 166322 76084
rect 171226 76032 171232 76084
rect 171284 76072 171290 76084
rect 171870 76072 171876 76084
rect 171284 76044 171876 76072
rect 171284 76032 171290 76044
rect 171870 76032 171876 76044
rect 171928 76032 171934 76084
rect 132862 75964 132868 76016
rect 132920 76004 132926 76016
rect 133874 76004 133880 76016
rect 132920 75976 133880 76004
rect 132920 75964 132926 75976
rect 133874 75964 133880 75976
rect 133932 75964 133938 76016
rect 134058 75964 134064 76016
rect 134116 76004 134122 76016
rect 134426 76004 134432 76016
rect 134116 75976 134432 76004
rect 134116 75964 134122 75976
rect 134426 75964 134432 75976
rect 134484 75964 134490 76016
rect 138474 75964 138480 76016
rect 138532 76004 138538 76016
rect 139118 76004 139124 76016
rect 138532 75976 139124 76004
rect 138532 75964 138538 75976
rect 139118 75964 139124 75976
rect 139176 75964 139182 76016
rect 151078 75964 151084 76016
rect 151136 76004 151142 76016
rect 151354 76004 151360 76016
rect 151136 75976 151360 76004
rect 151136 75964 151142 75976
rect 151354 75964 151360 75976
rect 151412 75964 151418 76016
rect 170674 75964 170680 76016
rect 170732 76004 170738 76016
rect 172054 76004 172060 76016
rect 170732 75976 172060 76004
rect 170732 75964 170738 75976
rect 172054 75964 172060 75976
rect 172112 75964 172118 76016
rect 130378 75896 130384 75948
rect 130436 75936 130442 75948
rect 154298 75936 154304 75948
rect 130436 75908 154304 75936
rect 130436 75896 130442 75908
rect 154298 75896 154304 75908
rect 154356 75896 154362 75948
rect 158990 75896 158996 75948
rect 159048 75936 159054 75948
rect 159266 75936 159272 75948
rect 159048 75908 159272 75936
rect 159048 75896 159054 75908
rect 159266 75896 159272 75908
rect 159324 75896 159330 75948
rect 159910 75896 159916 75948
rect 159968 75936 159974 75948
rect 160554 75936 160560 75948
rect 159968 75908 160560 75936
rect 159968 75896 159974 75908
rect 160554 75896 160560 75908
rect 160612 75896 160618 75948
rect 161750 75896 161756 75948
rect 161808 75936 161814 75948
rect 162118 75936 162124 75948
rect 161808 75908 162124 75936
rect 161808 75896 161814 75908
rect 162118 75896 162124 75908
rect 162176 75896 162182 75948
rect 168466 75896 168472 75948
rect 168524 75936 168530 75948
rect 168834 75936 168840 75948
rect 168524 75908 168840 75936
rect 168524 75896 168530 75908
rect 168834 75896 168840 75908
rect 168892 75896 168898 75948
rect 169938 75896 169944 75948
rect 169996 75936 170002 75948
rect 170122 75936 170128 75948
rect 169996 75908 170128 75936
rect 169996 75896 170002 75908
rect 170122 75896 170128 75908
rect 170180 75896 170186 75948
rect 171318 75896 171324 75948
rect 171376 75936 171382 75948
rect 171686 75936 171692 75948
rect 171376 75908 171692 75936
rect 171376 75896 171382 75908
rect 171686 75896 171692 75908
rect 171744 75896 171750 75948
rect 173342 75896 173348 75948
rect 173400 75936 173406 75948
rect 173710 75936 173716 75948
rect 173400 75908 173716 75936
rect 173400 75896 173406 75908
rect 173710 75896 173716 75908
rect 173768 75896 173774 75948
rect 176746 75896 176752 75948
rect 176804 75936 176810 75948
rect 177666 75936 177672 75948
rect 176804 75908 177672 75936
rect 176804 75896 176810 75908
rect 177666 75896 177672 75908
rect 177724 75896 177730 75948
rect 100386 75828 100392 75880
rect 100444 75868 100450 75880
rect 102134 75868 102140 75880
rect 100444 75840 102140 75868
rect 100444 75828 100450 75840
rect 102134 75828 102140 75840
rect 102192 75828 102198 75880
rect 150158 75868 150164 75880
rect 103486 75840 150164 75868
rect 97350 75760 97356 75812
rect 97408 75800 97414 75812
rect 103486 75800 103514 75840
rect 150158 75828 150164 75840
rect 150216 75828 150222 75880
rect 151078 75828 151084 75880
rect 151136 75868 151142 75880
rect 151630 75868 151636 75880
rect 151136 75840 151636 75868
rect 151136 75828 151142 75840
rect 151630 75828 151636 75840
rect 151688 75828 151694 75880
rect 160278 75828 160284 75880
rect 160336 75868 160342 75880
rect 160830 75868 160836 75880
rect 160336 75840 160836 75868
rect 160336 75828 160342 75840
rect 160830 75828 160836 75840
rect 160888 75828 160894 75880
rect 168742 75828 168748 75880
rect 168800 75868 168806 75880
rect 171778 75868 171784 75880
rect 168800 75840 171784 75868
rect 168800 75828 168806 75840
rect 171778 75828 171784 75840
rect 171836 75828 171842 75880
rect 172238 75828 172244 75880
rect 172296 75868 172302 75880
rect 191926 75868 191932 75880
rect 172296 75840 191932 75868
rect 172296 75828 172302 75840
rect 191926 75828 191932 75840
rect 191984 75828 191990 75880
rect 97408 75772 103514 75800
rect 97408 75760 97414 75772
rect 129642 75760 129648 75812
rect 129700 75800 129706 75812
rect 152826 75800 152832 75812
rect 129700 75772 152832 75800
rect 129700 75760 129706 75772
rect 152826 75760 152832 75772
rect 152884 75760 152890 75812
rect 169846 75760 169852 75812
rect 169904 75800 169910 75812
rect 170858 75800 170864 75812
rect 169904 75772 170864 75800
rect 169904 75760 169910 75772
rect 170858 75760 170864 75772
rect 170916 75760 170922 75812
rect 171594 75760 171600 75812
rect 171652 75800 171658 75812
rect 192938 75800 192944 75812
rect 171652 75772 192944 75800
rect 171652 75760 171658 75772
rect 192938 75760 192944 75772
rect 192996 75760 193002 75812
rect 117314 75692 117320 75744
rect 117372 75732 117378 75744
rect 121086 75732 121092 75744
rect 117372 75704 121092 75732
rect 117372 75692 117378 75704
rect 121086 75692 121092 75704
rect 121144 75732 121150 75744
rect 155770 75732 155776 75744
rect 121144 75704 155776 75732
rect 121144 75692 121150 75704
rect 155770 75692 155776 75704
rect 155828 75692 155834 75744
rect 175550 75692 175556 75744
rect 175608 75732 175614 75744
rect 215386 75732 215392 75744
rect 175608 75704 215392 75732
rect 175608 75692 175614 75704
rect 215386 75692 215392 75704
rect 215444 75732 215450 75744
rect 215846 75732 215852 75744
rect 215444 75704 215852 75732
rect 215444 75692 215450 75704
rect 215846 75692 215852 75704
rect 215904 75692 215910 75744
rect 117038 75624 117044 75676
rect 117096 75664 117102 75676
rect 149238 75664 149244 75676
rect 117096 75636 149244 75664
rect 117096 75624 117102 75636
rect 149238 75624 149244 75636
rect 149296 75664 149302 75676
rect 150158 75664 150164 75676
rect 149296 75636 150164 75664
rect 149296 75624 149302 75636
rect 150158 75624 150164 75636
rect 150216 75624 150222 75676
rect 175826 75624 175832 75676
rect 175884 75664 175890 75676
rect 215478 75664 215484 75676
rect 175884 75636 215484 75664
rect 175884 75624 175890 75636
rect 215478 75624 215484 75636
rect 215536 75624 215542 75676
rect 112806 75556 112812 75608
rect 112864 75596 112870 75608
rect 145926 75596 145932 75608
rect 112864 75568 145932 75596
rect 112864 75556 112870 75568
rect 145926 75556 145932 75568
rect 145984 75556 145990 75608
rect 170766 75556 170772 75608
rect 170824 75596 170830 75608
rect 208486 75596 208492 75608
rect 170824 75568 208492 75596
rect 170824 75556 170830 75568
rect 208486 75556 208492 75568
rect 208544 75556 208550 75608
rect 103238 75488 103244 75540
rect 103296 75528 103302 75540
rect 135254 75528 135260 75540
rect 103296 75500 135260 75528
rect 103296 75488 103302 75500
rect 36538 75216 36544 75268
rect 36596 75256 36602 75268
rect 103486 75256 103514 75500
rect 135254 75488 135260 75500
rect 135312 75488 135318 75540
rect 146662 75528 146668 75540
rect 140056 75500 146668 75528
rect 114370 75420 114376 75472
rect 114428 75460 114434 75472
rect 139946 75460 139952 75472
rect 114428 75432 139952 75460
rect 114428 75420 114434 75432
rect 139946 75420 139952 75432
rect 140004 75420 140010 75472
rect 116946 75352 116952 75404
rect 117004 75392 117010 75404
rect 140056 75392 140084 75500
rect 146662 75488 146668 75500
rect 146720 75488 146726 75540
rect 158254 75488 158260 75540
rect 158312 75528 158318 75540
rect 160646 75528 160652 75540
rect 158312 75500 160652 75528
rect 158312 75488 158318 75500
rect 160646 75488 160652 75500
rect 160704 75528 160710 75540
rect 195146 75528 195152 75540
rect 160704 75500 195152 75528
rect 160704 75488 160710 75500
rect 195146 75488 195152 75500
rect 195204 75488 195210 75540
rect 142246 75420 142252 75472
rect 142304 75460 142310 75472
rect 146202 75460 146208 75472
rect 142304 75432 146208 75460
rect 142304 75420 142310 75432
rect 146202 75420 146208 75432
rect 146260 75420 146266 75472
rect 156046 75420 156052 75472
rect 156104 75460 156110 75472
rect 157058 75460 157064 75472
rect 156104 75432 157064 75460
rect 156104 75420 156110 75432
rect 157058 75420 157064 75432
rect 157116 75420 157122 75472
rect 174538 75420 174544 75472
rect 174596 75460 174602 75472
rect 208578 75460 208584 75472
rect 174596 75432 208584 75460
rect 174596 75420 174602 75432
rect 208578 75420 208584 75432
rect 208636 75420 208642 75472
rect 145098 75392 145104 75404
rect 117004 75364 140084 75392
rect 140792 75364 145104 75392
rect 117004 75352 117010 75364
rect 117866 75284 117872 75336
rect 117924 75324 117930 75336
rect 140792 75324 140820 75364
rect 145098 75352 145104 75364
rect 145156 75352 145162 75404
rect 146386 75352 146392 75404
rect 146444 75392 146450 75404
rect 146846 75392 146852 75404
rect 146444 75364 146852 75392
rect 146444 75352 146450 75364
rect 146846 75352 146852 75364
rect 146904 75352 146910 75404
rect 157306 75364 166994 75392
rect 117924 75296 140820 75324
rect 117924 75284 117930 75296
rect 140866 75284 140872 75336
rect 140924 75324 140930 75336
rect 141970 75324 141976 75336
rect 140924 75296 141976 75324
rect 140924 75284 140930 75296
rect 141970 75284 141976 75296
rect 142028 75284 142034 75336
rect 142338 75284 142344 75336
rect 142396 75324 142402 75336
rect 142890 75324 142896 75336
rect 142396 75296 142896 75324
rect 142396 75284 142402 75296
rect 142890 75284 142896 75296
rect 142948 75284 142954 75336
rect 142982 75284 142988 75336
rect 143040 75324 143046 75336
rect 143040 75296 147674 75324
rect 143040 75284 143046 75296
rect 36596 75228 103514 75256
rect 36596 75216 36602 75228
rect 134242 75216 134248 75268
rect 134300 75256 134306 75268
rect 134794 75256 134800 75268
rect 134300 75228 134800 75256
rect 134300 75216 134306 75228
rect 134794 75216 134800 75228
rect 134852 75216 134858 75268
rect 137002 75216 137008 75268
rect 137060 75256 137066 75268
rect 137646 75256 137652 75268
rect 137060 75228 137652 75256
rect 137060 75216 137066 75228
rect 137646 75216 137652 75228
rect 137704 75216 137710 75268
rect 139946 75216 139952 75268
rect 140004 75256 140010 75268
rect 142246 75256 142252 75268
rect 140004 75228 142252 75256
rect 140004 75216 140010 75228
rect 142246 75216 142252 75228
rect 142304 75216 142310 75268
rect 142614 75216 142620 75268
rect 142672 75256 142678 75268
rect 142798 75256 142804 75268
rect 142672 75228 142804 75256
rect 142672 75216 142678 75228
rect 142798 75216 142804 75228
rect 142856 75216 142862 75268
rect 143902 75216 143908 75268
rect 143960 75256 143966 75268
rect 144270 75256 144276 75268
rect 143960 75228 144276 75256
rect 143960 75216 143966 75228
rect 144270 75216 144276 75228
rect 144328 75216 144334 75268
rect 147646 75256 147674 75296
rect 157306 75256 157334 75364
rect 147646 75228 157334 75256
rect 164234 75216 164240 75268
rect 164292 75256 164298 75268
rect 164602 75256 164608 75268
rect 164292 75228 164608 75256
rect 164292 75216 164298 75228
rect 164602 75216 164608 75228
rect 164660 75216 164666 75268
rect 78674 75148 78680 75200
rect 78732 75188 78738 75200
rect 78732 75160 147674 75188
rect 78732 75148 78738 75160
rect 108850 75080 108856 75132
rect 108908 75120 108914 75132
rect 108908 75092 138014 75120
rect 108908 75080 108914 75092
rect 108482 75012 108488 75064
rect 108540 75052 108546 75064
rect 132126 75052 132132 75064
rect 108540 75024 132132 75052
rect 108540 75012 108546 75024
rect 132126 75012 132132 75024
rect 132184 75012 132190 75064
rect 134150 75012 134156 75064
rect 134208 75052 134214 75064
rect 134518 75052 134524 75064
rect 134208 75024 134524 75052
rect 134208 75012 134214 75024
rect 134518 75012 134524 75024
rect 134576 75012 134582 75064
rect 137986 75052 138014 75092
rect 141050 75080 141056 75132
rect 141108 75120 141114 75132
rect 141878 75120 141884 75132
rect 141108 75092 141884 75120
rect 141108 75080 141114 75092
rect 141878 75080 141884 75092
rect 141936 75080 141942 75132
rect 142522 75052 142528 75064
rect 137986 75024 142528 75052
rect 142522 75012 142528 75024
rect 142580 75052 142586 75064
rect 142982 75052 142988 75064
rect 142580 75024 142988 75052
rect 142580 75012 142586 75024
rect 142982 75012 142988 75024
rect 143040 75012 143046 75064
rect 147646 75052 147674 75160
rect 148134 75148 148140 75200
rect 148192 75188 148198 75200
rect 148318 75188 148324 75200
rect 148192 75160 148324 75188
rect 148192 75148 148198 75160
rect 148318 75148 148324 75160
rect 148376 75148 148382 75200
rect 164326 75148 164332 75200
rect 164384 75188 164390 75200
rect 165338 75188 165344 75200
rect 164384 75160 165344 75188
rect 164384 75148 164390 75160
rect 165338 75148 165344 75160
rect 165396 75148 165402 75200
rect 163406 75080 163412 75132
rect 163464 75120 163470 75132
rect 166966 75120 166994 75364
rect 169202 75352 169208 75404
rect 169260 75392 169266 75404
rect 201770 75392 201776 75404
rect 169260 75364 201776 75392
rect 169260 75352 169266 75364
rect 201770 75352 201776 75364
rect 201828 75392 201834 75404
rect 202782 75392 202788 75404
rect 201828 75364 202788 75392
rect 201828 75352 201834 75364
rect 202782 75352 202788 75364
rect 202840 75352 202846 75404
rect 180518 75284 180524 75336
rect 180576 75324 180582 75336
rect 210234 75324 210240 75336
rect 180576 75296 210240 75324
rect 180576 75284 180582 75296
rect 210234 75284 210240 75296
rect 210292 75284 210298 75336
rect 167178 75216 167184 75268
rect 167236 75256 167242 75268
rect 167730 75256 167736 75268
rect 167236 75228 167736 75256
rect 167236 75216 167242 75228
rect 167730 75216 167736 75228
rect 167788 75216 167794 75268
rect 174078 75216 174084 75268
rect 174136 75256 174142 75268
rect 174354 75256 174360 75268
rect 174136 75228 174360 75256
rect 174136 75216 174142 75228
rect 174354 75216 174360 75228
rect 174412 75216 174418 75268
rect 202782 75216 202788 75268
rect 202840 75256 202846 75268
rect 281534 75256 281540 75268
rect 202840 75228 281540 75256
rect 202840 75216 202846 75228
rect 281534 75216 281540 75228
rect 281592 75216 281598 75268
rect 167086 75148 167092 75200
rect 167144 75188 167150 75200
rect 168282 75188 168288 75200
rect 167144 75160 168288 75188
rect 167144 75148 167150 75160
rect 168282 75148 168288 75160
rect 168340 75148 168346 75200
rect 181438 75148 181444 75200
rect 181496 75188 181502 75200
rect 214098 75188 214104 75200
rect 181496 75160 214104 75188
rect 181496 75148 181502 75160
rect 214098 75148 214104 75160
rect 214156 75148 214162 75200
rect 215386 75148 215392 75200
rect 215444 75188 215450 75200
rect 525794 75188 525800 75200
rect 215444 75160 525800 75188
rect 215444 75148 215450 75160
rect 525794 75148 525800 75160
rect 525852 75148 525858 75200
rect 174538 75120 174544 75132
rect 163464 75092 165752 75120
rect 166966 75092 174544 75120
rect 163464 75080 163470 75092
rect 158254 75052 158260 75064
rect 147646 75024 158260 75052
rect 158254 75012 158260 75024
rect 158312 75012 158318 75064
rect 164234 75012 164240 75064
rect 164292 75052 164298 75064
rect 165154 75052 165160 75064
rect 164292 75024 165160 75052
rect 164292 75012 164298 75024
rect 165154 75012 165160 75024
rect 165212 75012 165218 75064
rect 165724 75052 165752 75092
rect 174538 75080 174544 75092
rect 174596 75080 174602 75132
rect 177942 75080 177948 75132
rect 178000 75120 178006 75132
rect 207290 75120 207296 75132
rect 178000 75092 207296 75120
rect 178000 75080 178006 75092
rect 207290 75080 207296 75092
rect 207348 75080 207354 75132
rect 214650 75052 214656 75064
rect 165724 75024 214656 75052
rect 214650 75012 214656 75024
rect 214708 75012 214714 75064
rect 120350 74944 120356 74996
rect 120408 74984 120414 74996
rect 142430 74984 142436 74996
rect 120408 74956 142436 74984
rect 120408 74944 120414 74956
rect 142430 74944 142436 74956
rect 142488 74984 142494 74996
rect 142798 74984 142804 74996
rect 142488 74956 142804 74984
rect 142488 74944 142494 74956
rect 142798 74944 142804 74956
rect 142856 74944 142862 74996
rect 157150 74944 157156 74996
rect 157208 74984 157214 74996
rect 214742 74984 214748 74996
rect 157208 74956 214748 74984
rect 157208 74944 157214 74956
rect 214742 74944 214748 74956
rect 214800 74944 214806 74996
rect 149698 74876 149704 74928
rect 149756 74916 149762 74928
rect 179966 74916 179972 74928
rect 149756 74888 179972 74916
rect 149756 74876 149762 74888
rect 179966 74876 179972 74888
rect 180024 74876 180030 74928
rect 161290 74808 161296 74860
rect 161348 74848 161354 74860
rect 181806 74848 181812 74860
rect 161348 74820 181812 74848
rect 161348 74808 161354 74820
rect 181806 74808 181812 74820
rect 181864 74808 181870 74860
rect 167178 74740 167184 74792
rect 167236 74780 167242 74792
rect 168098 74780 168104 74792
rect 167236 74752 168104 74780
rect 167236 74740 167242 74752
rect 168098 74740 168104 74752
rect 168156 74740 168162 74792
rect 153930 74604 153936 74656
rect 153988 74644 153994 74656
rect 154206 74644 154212 74656
rect 153988 74616 154212 74644
rect 153988 74604 153994 74616
rect 154206 74604 154212 74616
rect 154264 74604 154270 74656
rect 107286 74468 107292 74520
rect 107344 74508 107350 74520
rect 132402 74508 132408 74520
rect 107344 74480 132408 74508
rect 107344 74468 107350 74480
rect 132402 74468 132408 74480
rect 132460 74468 132466 74520
rect 169294 74468 169300 74520
rect 169352 74508 169358 74520
rect 191006 74508 191012 74520
rect 169352 74480 191012 74508
rect 169352 74468 169358 74480
rect 191006 74468 191012 74480
rect 191064 74468 191070 74520
rect 127526 74400 127532 74452
rect 127584 74440 127590 74452
rect 147766 74440 147772 74452
rect 127584 74412 147772 74440
rect 127584 74400 127590 74412
rect 147766 74400 147772 74412
rect 147824 74400 147830 74452
rect 175734 74400 175740 74452
rect 175792 74440 175798 74452
rect 211706 74440 211712 74452
rect 175792 74412 211712 74440
rect 175792 74400 175798 74412
rect 211706 74400 211712 74412
rect 211764 74400 211770 74452
rect 120534 74332 120540 74384
rect 120592 74372 120598 74384
rect 158622 74372 158628 74384
rect 120592 74344 158628 74372
rect 120592 74332 120598 74344
rect 158622 74332 158628 74344
rect 158680 74332 158686 74384
rect 162302 74332 162308 74384
rect 162360 74372 162366 74384
rect 196526 74372 196532 74384
rect 162360 74344 196532 74372
rect 162360 74332 162366 74344
rect 196526 74332 196532 74344
rect 196584 74332 196590 74384
rect 109770 74264 109776 74316
rect 109828 74304 109834 74316
rect 143534 74304 143540 74316
rect 109828 74276 143540 74304
rect 109828 74264 109834 74276
rect 143534 74264 143540 74276
rect 143592 74264 143598 74316
rect 159450 74264 159456 74316
rect 159508 74304 159514 74316
rect 192294 74304 192300 74316
rect 159508 74276 192300 74304
rect 159508 74264 159514 74276
rect 192294 74264 192300 74276
rect 192352 74264 192358 74316
rect 114738 74196 114744 74248
rect 114796 74236 114802 74248
rect 147674 74236 147680 74248
rect 114796 74208 147680 74236
rect 114796 74196 114802 74208
rect 147674 74196 147680 74208
rect 147732 74196 147738 74248
rect 166626 74196 166632 74248
rect 166684 74236 166690 74248
rect 197446 74236 197452 74248
rect 166684 74208 197452 74236
rect 166684 74196 166690 74208
rect 197446 74196 197452 74208
rect 197504 74196 197510 74248
rect 119982 74128 119988 74180
rect 120040 74168 120046 74180
rect 152366 74168 152372 74180
rect 120040 74140 152372 74168
rect 120040 74128 120046 74140
rect 152366 74128 152372 74140
rect 152424 74128 152430 74180
rect 165614 74128 165620 74180
rect 165672 74168 165678 74180
rect 196158 74168 196164 74180
rect 165672 74140 196164 74168
rect 165672 74128 165678 74140
rect 196158 74128 196164 74140
rect 196216 74128 196222 74180
rect 113910 74060 113916 74112
rect 113968 74100 113974 74112
rect 145742 74100 145748 74112
rect 113968 74072 145748 74100
rect 113968 74060 113974 74072
rect 145742 74060 145748 74072
rect 145800 74060 145806 74112
rect 163866 74060 163872 74112
rect 163924 74100 163930 74112
rect 193858 74100 193864 74112
rect 163924 74072 193864 74100
rect 163924 74060 163930 74072
rect 193858 74060 193864 74072
rect 193916 74060 193922 74112
rect 119522 73992 119528 74044
rect 119580 74032 119586 74044
rect 151446 74032 151452 74044
rect 119580 74004 151452 74032
rect 119580 73992 119586 74004
rect 151446 73992 151452 74004
rect 151504 73992 151510 74044
rect 159726 73992 159732 74044
rect 159784 74032 159790 74044
rect 193582 74032 193588 74044
rect 159784 74004 193588 74032
rect 159784 73992 159790 74004
rect 193582 73992 193588 74004
rect 193640 73992 193646 74044
rect 115382 73924 115388 73976
rect 115440 73964 115446 73976
rect 145282 73964 145288 73976
rect 115440 73936 145288 73964
rect 115440 73924 115446 73936
rect 145282 73924 145288 73936
rect 145340 73924 145346 73976
rect 172514 73924 172520 73976
rect 172572 73964 172578 73976
rect 199286 73964 199292 73976
rect 172572 73936 199292 73964
rect 172572 73924 172578 73936
rect 199286 73924 199292 73936
rect 199344 73924 199350 73976
rect 114002 73856 114008 73908
rect 114060 73896 114066 73908
rect 142154 73896 142160 73908
rect 114060 73868 142160 73896
rect 114060 73856 114066 73868
rect 142154 73856 142160 73868
rect 142212 73856 142218 73908
rect 162670 73856 162676 73908
rect 162728 73896 162734 73908
rect 182174 73896 182180 73908
rect 162728 73868 182180 73896
rect 162728 73856 162734 73868
rect 182174 73856 182180 73868
rect 182232 73856 182238 73908
rect 13078 73788 13084 73840
rect 13136 73828 13142 73840
rect 119522 73828 119528 73840
rect 13136 73800 119528 73828
rect 13136 73788 13142 73800
rect 119522 73788 119528 73800
rect 119580 73788 119586 73840
rect 143534 73788 143540 73840
rect 143592 73828 143598 73840
rect 144178 73828 144184 73840
rect 143592 73800 144184 73828
rect 143592 73788 143598 73800
rect 144178 73788 144184 73800
rect 144236 73828 144242 73840
rect 274634 73828 274640 73840
rect 144236 73800 274640 73828
rect 144236 73788 144242 73800
rect 274634 73788 274640 73800
rect 274692 73788 274698 73840
rect 107470 73720 107476 73772
rect 107528 73760 107534 73772
rect 132034 73760 132040 73772
rect 107528 73732 132040 73760
rect 107528 73720 107534 73732
rect 132034 73720 132040 73732
rect 132092 73720 132098 73772
rect 164694 73720 164700 73772
rect 164752 73760 164758 73772
rect 202966 73760 202972 73772
rect 164752 73732 202972 73760
rect 164752 73720 164758 73732
rect 202966 73720 202972 73732
rect 203024 73720 203030 73772
rect 94774 73652 94780 73704
rect 94832 73692 94838 73704
rect 148870 73692 148876 73704
rect 94832 73664 148876 73692
rect 94832 73652 94838 73664
rect 148870 73652 148876 73664
rect 148928 73652 148934 73704
rect 165982 73652 165988 73704
rect 166040 73692 166046 73704
rect 190730 73692 190736 73704
rect 166040 73664 190736 73692
rect 166040 73652 166046 73664
rect 190730 73652 190736 73664
rect 190788 73652 190794 73704
rect 109586 73584 109592 73636
rect 109644 73624 109650 73636
rect 148042 73624 148048 73636
rect 109644 73596 148048 73624
rect 109644 73584 109650 73596
rect 148042 73584 148048 73596
rect 148100 73584 148106 73636
rect 182082 73584 182088 73636
rect 182140 73624 182146 73636
rect 201678 73624 201684 73636
rect 182140 73596 201684 73624
rect 182140 73584 182146 73596
rect 201678 73584 201684 73596
rect 201736 73584 201742 73636
rect 105538 73516 105544 73568
rect 105596 73556 105602 73568
rect 131206 73556 131212 73568
rect 105596 73528 131212 73556
rect 105596 73516 105602 73528
rect 131206 73516 131212 73528
rect 131264 73516 131270 73568
rect 3142 73108 3148 73160
rect 3200 73148 3206 73160
rect 111794 73148 111800 73160
rect 3200 73120 111800 73148
rect 3200 73108 3206 73120
rect 111794 73108 111800 73120
rect 111852 73108 111858 73160
rect 123570 73108 123576 73160
rect 123628 73148 123634 73160
rect 123628 73120 128354 73148
rect 123628 73108 123634 73120
rect 128326 73080 128354 73120
rect 129274 73108 129280 73160
rect 129332 73148 129338 73160
rect 152090 73148 152096 73160
rect 129332 73120 152096 73148
rect 129332 73108 129338 73120
rect 152090 73108 152096 73120
rect 152148 73108 152154 73160
rect 158162 73108 158168 73160
rect 158220 73148 158226 73160
rect 158622 73148 158628 73160
rect 158220 73120 158628 73148
rect 158220 73108 158226 73120
rect 158622 73108 158628 73120
rect 158680 73108 158686 73160
rect 182174 73108 182180 73160
rect 182232 73148 182238 73160
rect 183462 73148 183468 73160
rect 182232 73120 183468 73148
rect 182232 73108 182238 73120
rect 183462 73108 183468 73120
rect 183520 73148 183526 73160
rect 193674 73148 193680 73160
rect 183520 73120 193680 73148
rect 183520 73108 183526 73120
rect 193674 73108 193680 73120
rect 193732 73108 193738 73160
rect 131206 73080 131212 73092
rect 128326 73052 131212 73080
rect 131206 73040 131212 73052
rect 131264 73080 131270 73092
rect 132310 73080 132316 73092
rect 131264 73052 132316 73080
rect 131264 73040 131270 73052
rect 132310 73040 132316 73052
rect 132368 73040 132374 73092
rect 138934 73040 138940 73092
rect 138992 73080 138998 73092
rect 143626 73080 143632 73092
rect 138992 73052 143632 73080
rect 138992 73040 138998 73052
rect 143626 73040 143632 73052
rect 143684 73040 143690 73092
rect 144086 73040 144092 73092
rect 144144 73080 144150 73092
rect 144454 73080 144460 73092
rect 144144 73052 144460 73080
rect 144144 73040 144150 73052
rect 144454 73040 144460 73052
rect 144512 73040 144518 73092
rect 172330 73040 172336 73092
rect 172388 73080 172394 73092
rect 203794 73080 203800 73092
rect 172388 73052 203800 73080
rect 172388 73040 172394 73052
rect 203794 73040 203800 73052
rect 203852 73040 203858 73092
rect 112714 72972 112720 73024
rect 112772 73012 112778 73024
rect 138750 73012 138756 73024
rect 112772 72984 138756 73012
rect 112772 72972 112778 72984
rect 138750 72972 138756 72984
rect 138808 72972 138814 73024
rect 142982 72972 142988 73024
rect 143040 73012 143046 73024
rect 143166 73012 143172 73024
rect 143040 72984 143172 73012
rect 143040 72972 143046 72984
rect 143166 72972 143172 72984
rect 143224 72972 143230 73024
rect 166258 72972 166264 73024
rect 166316 73012 166322 73024
rect 196710 73012 196716 73024
rect 166316 72984 196716 73012
rect 166316 72972 166322 72984
rect 196710 72972 196716 72984
rect 196768 72972 196774 73024
rect 126330 72904 126336 72956
rect 126388 72944 126394 72956
rect 150802 72944 150808 72956
rect 126388 72916 150808 72944
rect 126388 72904 126394 72916
rect 150802 72904 150808 72916
rect 150860 72904 150866 72956
rect 156782 72904 156788 72956
rect 156840 72944 156846 72956
rect 190914 72944 190920 72956
rect 156840 72916 190920 72944
rect 156840 72904 156846 72916
rect 190914 72904 190920 72916
rect 190972 72944 190978 72956
rect 191742 72944 191748 72956
rect 190972 72916 191748 72944
rect 190972 72904 190978 72916
rect 191742 72904 191748 72916
rect 191800 72904 191806 72956
rect 101950 72836 101956 72888
rect 102008 72876 102014 72888
rect 106274 72876 106280 72888
rect 102008 72848 106280 72876
rect 102008 72836 102014 72848
rect 106274 72836 106280 72848
rect 106332 72876 106338 72888
rect 107470 72876 107476 72888
rect 106332 72848 107476 72876
rect 106332 72836 106338 72848
rect 107470 72836 107476 72848
rect 107528 72836 107534 72888
rect 118510 72836 118516 72888
rect 118568 72876 118574 72888
rect 151906 72876 151912 72888
rect 118568 72848 151912 72876
rect 118568 72836 118574 72848
rect 151906 72836 151912 72848
rect 151964 72836 151970 72888
rect 162578 72836 162584 72888
rect 162636 72876 162642 72888
rect 194686 72876 194692 72888
rect 162636 72848 194692 72876
rect 162636 72836 162642 72848
rect 194686 72836 194692 72848
rect 194744 72836 194750 72888
rect 119062 72768 119068 72820
rect 119120 72808 119126 72820
rect 153286 72808 153292 72820
rect 119120 72780 153292 72808
rect 119120 72768 119126 72780
rect 153286 72768 153292 72780
rect 153344 72768 153350 72820
rect 162762 72768 162768 72820
rect 162820 72808 162826 72820
rect 195974 72808 195980 72820
rect 162820 72780 195980 72808
rect 162820 72768 162826 72780
rect 195974 72768 195980 72780
rect 196032 72768 196038 72820
rect 113450 72700 113456 72752
rect 113508 72740 113514 72752
rect 147858 72740 147864 72752
rect 113508 72712 147864 72740
rect 113508 72700 113514 72712
rect 147858 72700 147864 72712
rect 147916 72700 147922 72752
rect 156506 72700 156512 72752
rect 156564 72740 156570 72752
rect 156782 72740 156788 72752
rect 156564 72712 156788 72740
rect 156564 72700 156570 72712
rect 156782 72700 156788 72712
rect 156840 72740 156846 72752
rect 190454 72740 190460 72752
rect 156840 72712 190460 72740
rect 156840 72700 156846 72712
rect 190454 72700 190460 72712
rect 190512 72700 190518 72752
rect 111518 72632 111524 72684
rect 111576 72672 111582 72684
rect 144454 72672 144460 72684
rect 111576 72644 144460 72672
rect 111576 72632 111582 72644
rect 144454 72632 144460 72644
rect 144512 72632 144518 72684
rect 158346 72632 158352 72684
rect 158404 72672 158410 72684
rect 189350 72672 189356 72684
rect 158404 72644 189356 72672
rect 158404 72632 158410 72644
rect 189350 72632 189356 72644
rect 189408 72632 189414 72684
rect 110230 72564 110236 72616
rect 110288 72604 110294 72616
rect 142982 72604 142988 72616
rect 110288 72576 142988 72604
rect 110288 72564 110294 72576
rect 142982 72564 142988 72576
rect 143040 72564 143046 72616
rect 175642 72564 175648 72616
rect 175700 72604 175706 72616
rect 204438 72604 204444 72616
rect 175700 72576 204444 72604
rect 175700 72564 175706 72576
rect 204438 72564 204444 72576
rect 204496 72564 204502 72616
rect 119706 72496 119712 72548
rect 119764 72536 119770 72548
rect 151814 72536 151820 72548
rect 119764 72508 151820 72536
rect 119764 72496 119770 72508
rect 151814 72496 151820 72508
rect 151872 72496 151878 72548
rect 169478 72496 169484 72548
rect 169536 72536 169542 72548
rect 194594 72536 194600 72548
rect 169536 72508 194600 72536
rect 169536 72496 169542 72508
rect 194594 72496 194600 72508
rect 194652 72496 194658 72548
rect 54478 72428 54484 72480
rect 54536 72468 54542 72480
rect 100294 72468 100300 72480
rect 54536 72440 100300 72468
rect 54536 72428 54542 72440
rect 100294 72428 100300 72440
rect 100352 72468 100358 72480
rect 134978 72468 134984 72480
rect 100352 72440 134984 72468
rect 100352 72428 100358 72440
rect 134978 72428 134984 72440
rect 135036 72428 135042 72480
rect 145190 72428 145196 72480
rect 145248 72468 145254 72480
rect 185578 72468 185584 72480
rect 145248 72440 185584 72468
rect 145248 72428 145254 72440
rect 185578 72428 185584 72440
rect 185636 72428 185642 72480
rect 191742 72428 191748 72480
rect 191800 72468 191806 72480
rect 255314 72468 255320 72480
rect 191800 72440 255320 72468
rect 191800 72428 191806 72440
rect 255314 72428 255320 72440
rect 255372 72428 255378 72480
rect 98638 72360 98644 72412
rect 98696 72400 98702 72412
rect 133782 72400 133788 72412
rect 98696 72372 133788 72400
rect 98696 72360 98702 72372
rect 133782 72360 133788 72372
rect 133840 72360 133846 72412
rect 158622 72360 158628 72412
rect 158680 72400 158686 72412
rect 192386 72400 192392 72412
rect 158680 72372 192392 72400
rect 158680 72360 158686 72372
rect 192386 72360 192392 72372
rect 192444 72360 192450 72412
rect 111794 72292 111800 72344
rect 111852 72332 111858 72344
rect 112622 72332 112628 72344
rect 111852 72304 112628 72332
rect 111852 72292 111858 72304
rect 112622 72292 112628 72304
rect 112680 72332 112686 72344
rect 147490 72332 147496 72344
rect 112680 72304 147496 72332
rect 112680 72292 112686 72304
rect 147490 72292 147496 72304
rect 147548 72292 147554 72344
rect 153838 72292 153844 72344
rect 153896 72332 153902 72344
rect 218054 72332 218060 72344
rect 153896 72304 218060 72332
rect 153896 72292 153902 72304
rect 218054 72292 218060 72304
rect 218112 72292 218118 72344
rect 94590 72224 94596 72276
rect 94648 72264 94654 72276
rect 157610 72264 157616 72276
rect 94648 72236 157616 72264
rect 94648 72224 94654 72236
rect 157610 72224 157616 72236
rect 157668 72224 157674 72276
rect 153930 72020 153936 72072
rect 153988 72060 153994 72072
rect 154206 72060 154212 72072
rect 153988 72032 154212 72060
rect 153988 72020 153994 72032
rect 154206 72020 154212 72032
rect 154264 72020 154270 72072
rect 108574 71680 108580 71732
rect 108632 71720 108638 71732
rect 143350 71720 143356 71732
rect 108632 71692 143356 71720
rect 108632 71680 108638 71692
rect 143350 71680 143356 71692
rect 143408 71680 143414 71732
rect 143718 71680 143724 71732
rect 143776 71720 143782 71732
rect 144178 71720 144184 71732
rect 143776 71692 144184 71720
rect 143776 71680 143782 71692
rect 144178 71680 144184 71692
rect 144236 71680 144242 71732
rect 173802 71680 173808 71732
rect 173860 71720 173866 71732
rect 174906 71720 174912 71732
rect 173860 71692 174912 71720
rect 173860 71680 173866 71692
rect 174906 71680 174912 71692
rect 174964 71680 174970 71732
rect 175274 71680 175280 71732
rect 175332 71720 175338 71732
rect 176102 71720 176108 71732
rect 175332 71692 176108 71720
rect 175332 71680 175338 71692
rect 176102 71680 176108 71692
rect 176160 71680 176166 71732
rect 210142 71720 210148 71732
rect 176212 71692 210148 71720
rect 114830 71612 114836 71664
rect 114888 71652 114894 71664
rect 149146 71652 149152 71664
rect 114888 71624 149152 71652
rect 114888 71612 114894 71624
rect 149146 71612 149152 71624
rect 149204 71652 149210 71664
rect 149882 71652 149888 71664
rect 149204 71624 149888 71652
rect 149204 71612 149210 71624
rect 149882 71612 149888 71624
rect 149940 71612 149946 71664
rect 169386 71612 169392 71664
rect 169444 71652 169450 71664
rect 176212 71652 176240 71692
rect 210142 71680 210148 71692
rect 210200 71680 210206 71732
rect 169444 71624 176240 71652
rect 169444 71612 169450 71624
rect 176562 71612 176568 71664
rect 176620 71652 176626 71664
rect 215294 71652 215300 71664
rect 176620 71624 215300 71652
rect 176620 71612 176626 71624
rect 215294 71612 215300 71624
rect 215352 71612 215358 71664
rect 119890 71544 119896 71596
rect 119948 71584 119954 71596
rect 153838 71584 153844 71596
rect 119948 71556 153844 71584
rect 119948 71544 119954 71556
rect 153838 71544 153844 71556
rect 153896 71544 153902 71596
rect 171410 71544 171416 71596
rect 171468 71584 171474 71596
rect 206002 71584 206008 71596
rect 171468 71556 206008 71584
rect 171468 71544 171474 71556
rect 206002 71544 206008 71556
rect 206060 71544 206066 71596
rect 207106 71544 207112 71596
rect 207164 71584 207170 71596
rect 207290 71584 207296 71596
rect 207164 71556 207296 71584
rect 207164 71544 207170 71556
rect 207290 71544 207296 71556
rect 207348 71544 207354 71596
rect 126238 71476 126244 71528
rect 126296 71516 126302 71528
rect 151078 71516 151084 71528
rect 126296 71488 151084 71516
rect 126296 71476 126302 71488
rect 151078 71476 151084 71488
rect 151136 71476 151142 71528
rect 170490 71476 170496 71528
rect 170548 71516 170554 71528
rect 204254 71516 204260 71528
rect 170548 71488 204260 71516
rect 170548 71476 170554 71488
rect 204254 71476 204260 71488
rect 204312 71476 204318 71528
rect 116670 71408 116676 71460
rect 116728 71448 116734 71460
rect 149790 71448 149796 71460
rect 116728 71420 149796 71448
rect 116728 71408 116734 71420
rect 149790 71408 149796 71420
rect 149848 71408 149854 71460
rect 165430 71408 165436 71460
rect 165488 71448 165494 71460
rect 197906 71448 197912 71460
rect 165488 71420 197912 71448
rect 165488 71408 165494 71420
rect 197906 71408 197912 71420
rect 197964 71408 197970 71460
rect 110782 71340 110788 71392
rect 110840 71380 110846 71392
rect 143718 71380 143724 71392
rect 110840 71352 143724 71380
rect 110840 71340 110846 71352
rect 143718 71340 143724 71352
rect 143776 71340 143782 71392
rect 174722 71340 174728 71392
rect 174780 71380 174786 71392
rect 207106 71380 207112 71392
rect 174780 71352 207112 71380
rect 174780 71340 174786 71352
rect 207106 71340 207112 71352
rect 207164 71340 207170 71392
rect 110966 71272 110972 71324
rect 111024 71312 111030 71324
rect 143534 71312 143540 71324
rect 111024 71284 143540 71312
rect 111024 71272 111030 71284
rect 143534 71272 143540 71284
rect 143592 71312 143598 71324
rect 147030 71312 147036 71324
rect 143592 71284 147036 71312
rect 143592 71272 143598 71284
rect 147030 71272 147036 71284
rect 147088 71272 147094 71324
rect 171778 71272 171784 71324
rect 171836 71312 171842 71324
rect 203150 71312 203156 71324
rect 171836 71284 203156 71312
rect 171836 71272 171842 71284
rect 203150 71272 203156 71284
rect 203208 71272 203214 71324
rect 110690 71204 110696 71256
rect 110748 71244 110754 71256
rect 144362 71244 144368 71256
rect 110748 71216 144368 71244
rect 110748 71204 110754 71216
rect 144362 71204 144368 71216
rect 144420 71204 144426 71256
rect 173434 71204 173440 71256
rect 173492 71244 173498 71256
rect 201678 71244 201684 71256
rect 173492 71216 201684 71244
rect 173492 71204 173498 71216
rect 201678 71204 201684 71216
rect 201736 71244 201742 71256
rect 202138 71244 202144 71256
rect 201736 71216 202144 71244
rect 201736 71204 201742 71216
rect 202138 71204 202144 71216
rect 202196 71204 202202 71256
rect 117682 71136 117688 71188
rect 117740 71176 117746 71188
rect 149514 71176 149520 71188
rect 117740 71148 149520 71176
rect 117740 71136 117746 71148
rect 149514 71136 149520 71148
rect 149572 71136 149578 71188
rect 171502 71136 171508 71188
rect 171560 71176 171566 71188
rect 199746 71176 199752 71188
rect 171560 71148 199752 71176
rect 171560 71136 171566 71148
rect 199746 71136 199752 71148
rect 199804 71136 199810 71188
rect 133690 71068 133696 71120
rect 133748 71108 133754 71120
rect 265618 71108 265624 71120
rect 133748 71080 265624 71108
rect 133748 71068 133754 71080
rect 265618 71068 265624 71080
rect 265676 71068 265682 71120
rect 4798 71000 4804 71052
rect 4856 71040 4862 71052
rect 156782 71040 156788 71052
rect 4856 71012 156788 71040
rect 4856 71000 4862 71012
rect 156782 71000 156788 71012
rect 156840 71000 156846 71052
rect 164786 71000 164792 71052
rect 164844 71040 164850 71052
rect 165338 71040 165344 71052
rect 164844 71012 165344 71040
rect 164844 71000 164850 71012
rect 165338 71000 165344 71012
rect 165396 71000 165402 71052
rect 176102 71000 176108 71052
rect 176160 71040 176166 71052
rect 199562 71040 199568 71052
rect 176160 71012 199568 71040
rect 176160 71000 176166 71012
rect 199562 71000 199568 71012
rect 199620 71000 199626 71052
rect 215294 71000 215300 71052
rect 215352 71040 215358 71052
rect 484394 71040 484400 71052
rect 215352 71012 484400 71040
rect 215352 71000 215358 71012
rect 484394 71000 484400 71012
rect 484452 71000 484458 71052
rect 111426 70932 111432 70984
rect 111484 70972 111490 70984
rect 140590 70972 140596 70984
rect 111484 70944 140596 70972
rect 111484 70932 111490 70944
rect 140590 70932 140596 70944
rect 140648 70932 140654 70984
rect 177022 70932 177028 70984
rect 177080 70972 177086 70984
rect 196342 70972 196348 70984
rect 177080 70944 196348 70972
rect 177080 70932 177086 70944
rect 196342 70932 196348 70944
rect 196400 70932 196406 70984
rect 101766 70864 101772 70916
rect 101824 70904 101830 70916
rect 136542 70904 136548 70916
rect 101824 70876 136548 70904
rect 101824 70864 101830 70876
rect 136542 70864 136548 70876
rect 136600 70864 136606 70916
rect 156414 70864 156420 70916
rect 156472 70904 156478 70916
rect 187050 70904 187056 70916
rect 156472 70876 187056 70904
rect 156472 70864 156478 70876
rect 187050 70864 187056 70876
rect 187108 70864 187114 70916
rect 125594 70388 125600 70440
rect 125652 70428 125658 70440
rect 173802 70428 173808 70440
rect 125652 70400 173808 70428
rect 125652 70388 125658 70400
rect 173802 70388 173808 70400
rect 173860 70388 173866 70440
rect 111610 70320 111616 70372
rect 111668 70360 111674 70372
rect 145374 70360 145380 70372
rect 111668 70332 145380 70360
rect 111668 70320 111674 70332
rect 145374 70320 145380 70332
rect 145432 70360 145438 70372
rect 145558 70360 145564 70372
rect 145432 70332 145564 70360
rect 145432 70320 145438 70332
rect 145558 70320 145564 70332
rect 145616 70320 145622 70372
rect 172606 70320 172612 70372
rect 172664 70360 172670 70372
rect 193398 70360 193404 70372
rect 172664 70332 193404 70360
rect 172664 70320 172670 70332
rect 193398 70320 193404 70332
rect 193456 70320 193462 70372
rect 120718 70252 120724 70304
rect 120776 70292 120782 70304
rect 154666 70292 154672 70304
rect 120776 70264 154672 70292
rect 120776 70252 120782 70264
rect 154666 70252 154672 70264
rect 154724 70252 154730 70304
rect 165890 70252 165896 70304
rect 165948 70292 165954 70304
rect 207750 70292 207756 70304
rect 165948 70264 207756 70292
rect 165948 70252 165954 70264
rect 207750 70252 207756 70264
rect 207808 70252 207814 70304
rect 114278 70184 114284 70236
rect 114336 70224 114342 70236
rect 146846 70224 146852 70236
rect 114336 70196 146852 70224
rect 114336 70184 114342 70196
rect 146846 70184 146852 70196
rect 146904 70184 146910 70236
rect 176746 70184 176752 70236
rect 176804 70224 176810 70236
rect 212902 70224 212908 70236
rect 176804 70196 212908 70224
rect 176804 70184 176810 70196
rect 212902 70184 212908 70196
rect 212960 70184 212966 70236
rect 116762 70116 116768 70168
rect 116820 70156 116826 70168
rect 151354 70156 151360 70168
rect 116820 70128 151360 70156
rect 116820 70116 116826 70128
rect 151354 70116 151360 70128
rect 151412 70116 151418 70168
rect 166074 70116 166080 70168
rect 166132 70156 166138 70168
rect 200206 70156 200212 70168
rect 166132 70128 200212 70156
rect 166132 70116 166138 70128
rect 200206 70116 200212 70128
rect 200264 70116 200270 70168
rect 120626 70048 120632 70100
rect 120684 70088 120690 70100
rect 151998 70088 152004 70100
rect 120684 70060 152004 70088
rect 120684 70048 120690 70060
rect 151998 70048 152004 70060
rect 152056 70048 152062 70100
rect 172054 70048 172060 70100
rect 172112 70088 172118 70100
rect 205634 70088 205640 70100
rect 172112 70060 205640 70088
rect 172112 70048 172118 70060
rect 205634 70048 205640 70060
rect 205692 70048 205698 70100
rect 118234 69980 118240 70032
rect 118292 70020 118298 70032
rect 150710 70020 150716 70032
rect 118292 69992 150716 70020
rect 118292 69980 118298 69992
rect 150710 69980 150716 69992
rect 150768 69980 150774 70032
rect 174170 69980 174176 70032
rect 174228 70020 174234 70032
rect 207382 70020 207388 70032
rect 174228 69992 207388 70020
rect 174228 69980 174234 69992
rect 207382 69980 207388 69992
rect 207440 70020 207446 70032
rect 207658 70020 207664 70032
rect 207440 69992 207664 70020
rect 207440 69980 207446 69992
rect 207658 69980 207664 69992
rect 207716 69980 207722 70032
rect 115566 69912 115572 69964
rect 115624 69952 115630 69964
rect 148594 69952 148600 69964
rect 115624 69924 148600 69952
rect 115624 69912 115630 69924
rect 148594 69912 148600 69924
rect 148652 69912 148658 69964
rect 167822 69912 167828 69964
rect 167880 69952 167886 69964
rect 201494 69952 201500 69964
rect 167880 69924 201500 69952
rect 167880 69912 167886 69924
rect 201494 69912 201500 69924
rect 201552 69912 201558 69964
rect 112898 69844 112904 69896
rect 112956 69884 112962 69896
rect 145466 69884 145472 69896
rect 112956 69856 145472 69884
rect 112956 69844 112962 69856
rect 145466 69844 145472 69856
rect 145524 69844 145530 69896
rect 171962 69844 171968 69896
rect 172020 69884 172026 69896
rect 204254 69884 204260 69896
rect 172020 69856 204260 69884
rect 172020 69844 172026 69856
rect 204254 69844 204260 69856
rect 204312 69844 204318 69896
rect 115842 69776 115848 69828
rect 115900 69816 115906 69828
rect 148226 69816 148232 69828
rect 115900 69788 148232 69816
rect 115900 69776 115906 69788
rect 148226 69776 148232 69788
rect 148284 69776 148290 69828
rect 173342 69776 173348 69828
rect 173400 69816 173406 69828
rect 205634 69816 205640 69828
rect 173400 69788 205640 69816
rect 173400 69776 173406 69788
rect 205634 69776 205640 69788
rect 205692 69776 205698 69828
rect 64138 69708 64144 69760
rect 64196 69748 64202 69760
rect 98730 69748 98736 69760
rect 64196 69720 98736 69748
rect 64196 69708 64202 69720
rect 98730 69708 98736 69720
rect 98788 69748 98794 69760
rect 132954 69748 132960 69760
rect 98788 69720 132960 69748
rect 98788 69708 98794 69720
rect 132954 69708 132960 69720
rect 133012 69708 133018 69760
rect 142798 69708 142804 69760
rect 142856 69748 142862 69760
rect 300854 69748 300860 69760
rect 142856 69720 300860 69748
rect 142856 69708 142862 69720
rect 300854 69708 300860 69720
rect 300912 69708 300918 69760
rect 43438 69640 43444 69692
rect 43496 69680 43502 69692
rect 115658 69680 115664 69692
rect 43496 69652 115664 69680
rect 43496 69640 43502 69652
rect 115658 69640 115664 69652
rect 115716 69680 115722 69692
rect 115842 69680 115848 69692
rect 115716 69652 115848 69680
rect 115716 69640 115722 69652
rect 115842 69640 115848 69652
rect 115900 69640 115906 69692
rect 143442 69640 143448 69692
rect 143500 69680 143506 69692
rect 173894 69680 173900 69692
rect 143500 69652 173900 69680
rect 143500 69640 143506 69652
rect 173894 69640 173900 69652
rect 173952 69640 173958 69692
rect 176838 69640 176844 69692
rect 176896 69680 176902 69692
rect 207290 69680 207296 69692
rect 176896 69652 207296 69680
rect 176896 69640 176902 69652
rect 207290 69640 207296 69652
rect 207348 69640 207354 69692
rect 207382 69640 207388 69692
rect 207440 69680 207446 69692
rect 407114 69680 407120 69692
rect 207440 69652 407120 69680
rect 207440 69640 207446 69652
rect 407114 69640 407120 69652
rect 407172 69640 407178 69692
rect 109678 69572 109684 69624
rect 109736 69612 109742 69624
rect 137370 69612 137376 69624
rect 109736 69584 137376 69612
rect 109736 69572 109742 69584
rect 137370 69572 137376 69584
rect 137428 69572 137434 69624
rect 167638 69572 167644 69624
rect 167696 69612 167702 69624
rect 197814 69612 197820 69624
rect 167696 69584 197820 69612
rect 167696 69572 167702 69584
rect 197814 69572 197820 69584
rect 197872 69572 197878 69624
rect 99282 69504 99288 69556
rect 99340 69544 99346 69556
rect 132770 69544 132776 69556
rect 99340 69516 132776 69544
rect 99340 69504 99346 69516
rect 132770 69504 132776 69516
rect 132828 69504 132834 69556
rect 156598 69504 156604 69556
rect 156656 69544 156662 69556
rect 218330 69544 218336 69556
rect 156656 69516 218336 69544
rect 156656 69504 156662 69516
rect 218330 69504 218336 69516
rect 218388 69504 218394 69556
rect 166074 69028 166080 69080
rect 166132 69068 166138 69080
rect 166258 69068 166264 69080
rect 166132 69040 166264 69068
rect 166132 69028 166138 69040
rect 166258 69028 166264 69040
rect 166316 69028 166322 69080
rect 97902 68960 97908 69012
rect 97960 69000 97966 69012
rect 131114 69000 131120 69012
rect 97960 68972 131120 69000
rect 97960 68960 97966 68972
rect 131114 68960 131120 68972
rect 131172 68960 131178 69012
rect 152734 68960 152740 69012
rect 152792 69000 152798 69012
rect 216122 69000 216128 69012
rect 152792 68972 216128 69000
rect 152792 68960 152798 68972
rect 216122 68960 216128 68972
rect 216180 69000 216186 69012
rect 579982 69000 579988 69012
rect 216180 68972 579988 69000
rect 216180 68960 216186 68972
rect 579982 68960 579988 68972
rect 580040 68960 580046 69012
rect 3142 68892 3148 68944
rect 3200 68932 3206 68944
rect 111886 68932 111892 68944
rect 3200 68904 111892 68932
rect 3200 68892 3206 68904
rect 111886 68892 111892 68904
rect 111944 68892 111950 68944
rect 121730 68892 121736 68944
rect 121788 68932 121794 68944
rect 141234 68932 141240 68944
rect 121788 68904 141240 68932
rect 121788 68892 121794 68904
rect 141234 68892 141240 68904
rect 141292 68892 141298 68944
rect 160462 68892 160468 68944
rect 160520 68932 160526 68944
rect 182818 68932 182824 68944
rect 160520 68904 182824 68932
rect 160520 68892 160526 68904
rect 182818 68892 182824 68904
rect 182876 68892 182882 68944
rect 95050 68824 95056 68876
rect 95108 68864 95114 68876
rect 155310 68864 155316 68876
rect 95108 68836 155316 68864
rect 95108 68824 95114 68836
rect 155310 68824 155316 68836
rect 155368 68824 155374 68876
rect 171870 68824 171876 68876
rect 171928 68864 171934 68876
rect 196434 68864 196440 68876
rect 171928 68836 196440 68864
rect 171928 68824 171934 68836
rect 196434 68824 196440 68836
rect 196492 68824 196498 68876
rect 122190 68756 122196 68808
rect 122248 68796 122254 68808
rect 122834 68796 122840 68808
rect 122248 68768 122840 68796
rect 122248 68756 122254 68768
rect 122834 68756 122840 68768
rect 122892 68796 122898 68808
rect 146570 68796 146576 68808
rect 122892 68768 146576 68796
rect 122892 68756 122898 68768
rect 146570 68756 146576 68768
rect 146628 68756 146634 68808
rect 161382 68756 161388 68808
rect 161440 68796 161446 68808
rect 194870 68796 194876 68808
rect 161440 68768 194876 68796
rect 161440 68756 161446 68768
rect 194870 68756 194876 68768
rect 194928 68756 194934 68808
rect 104802 68688 104808 68740
rect 104860 68728 104866 68740
rect 138658 68728 138664 68740
rect 104860 68700 138664 68728
rect 104860 68688 104866 68700
rect 138658 68688 138664 68700
rect 138716 68688 138722 68740
rect 157518 68688 157524 68740
rect 157576 68728 157582 68740
rect 191834 68728 191840 68740
rect 157576 68700 191840 68728
rect 157576 68688 157582 68700
rect 191834 68688 191840 68700
rect 191892 68688 191898 68740
rect 105906 68620 105912 68672
rect 105964 68660 105970 68672
rect 139486 68660 139492 68672
rect 105964 68632 139492 68660
rect 105964 68620 105970 68632
rect 139486 68620 139492 68632
rect 139544 68620 139550 68672
rect 161934 68620 161940 68672
rect 161992 68660 161998 68672
rect 162762 68660 162768 68672
rect 161992 68632 162768 68660
rect 161992 68620 161998 68632
rect 162762 68620 162768 68632
rect 162820 68620 162826 68672
rect 193490 68660 193496 68672
rect 162872 68632 193496 68660
rect 101858 68552 101864 68604
rect 101916 68592 101922 68604
rect 136358 68592 136364 68604
rect 101916 68564 136364 68592
rect 101916 68552 101922 68564
rect 136358 68552 136364 68564
rect 136416 68552 136422 68604
rect 107010 68484 107016 68536
rect 107068 68524 107074 68536
rect 139854 68524 139860 68536
rect 107068 68496 139860 68524
rect 107068 68484 107074 68496
rect 139854 68484 139860 68496
rect 139912 68484 139918 68536
rect 160002 68484 160008 68536
rect 160060 68524 160066 68536
rect 162872 68524 162900 68632
rect 193490 68620 193496 68632
rect 193548 68620 193554 68672
rect 195514 68592 195520 68604
rect 160060 68496 162900 68524
rect 162964 68564 195520 68592
rect 160060 68484 160066 68496
rect 110138 68416 110144 68468
rect 110196 68456 110202 68468
rect 141418 68456 141424 68468
rect 110196 68428 141424 68456
rect 110196 68416 110202 68428
rect 141418 68416 141424 68428
rect 141476 68416 141482 68468
rect 161290 68416 161296 68468
rect 161348 68456 161354 68468
rect 162964 68456 162992 68564
rect 195514 68552 195520 68564
rect 195572 68552 195578 68604
rect 171962 68484 171968 68536
rect 172020 68524 172026 68536
rect 196894 68524 196900 68536
rect 172020 68496 196900 68524
rect 172020 68484 172026 68496
rect 196894 68484 196900 68496
rect 196952 68484 196958 68536
rect 193766 68456 193772 68468
rect 161348 68428 162992 68456
rect 171888 68428 193772 68456
rect 161348 68416 161354 68428
rect 107194 68348 107200 68400
rect 107252 68388 107258 68400
rect 135622 68388 135628 68400
rect 107252 68360 135628 68388
rect 107252 68348 107258 68360
rect 135622 68348 135628 68360
rect 135680 68348 135686 68400
rect 159174 68348 159180 68400
rect 159232 68388 159238 68400
rect 171888 68388 171916 68428
rect 193766 68416 193772 68428
rect 193824 68416 193830 68468
rect 159232 68360 171916 68388
rect 159232 68348 159238 68360
rect 172054 68348 172060 68400
rect 172112 68388 172118 68400
rect 199654 68388 199660 68400
rect 172112 68360 199660 68388
rect 172112 68348 172118 68360
rect 199654 68348 199660 68360
rect 199712 68348 199718 68400
rect 134610 68280 134616 68332
rect 134668 68320 134674 68332
rect 211798 68320 211804 68332
rect 134668 68292 211804 68320
rect 134668 68280 134674 68292
rect 211798 68280 211804 68292
rect 211856 68280 211862 68332
rect 111702 68212 111708 68264
rect 111760 68252 111766 68264
rect 152550 68252 152556 68264
rect 111760 68224 152556 68252
rect 111760 68212 111766 68224
rect 152550 68212 152556 68224
rect 152608 68212 152614 68264
rect 168926 68212 168932 68264
rect 168984 68252 168990 68264
rect 190454 68252 190460 68264
rect 168984 68224 190460 68252
rect 168984 68212 168990 68224
rect 190454 68212 190460 68224
rect 190512 68252 190518 68264
rect 203610 68252 203616 68264
rect 190512 68224 203616 68252
rect 190512 68212 190518 68224
rect 203610 68212 203616 68224
rect 203668 68212 203674 68264
rect 111886 68144 111892 68196
rect 111944 68184 111950 68196
rect 113082 68184 113088 68196
rect 111944 68156 113088 68184
rect 111944 68144 111950 68156
rect 113082 68144 113088 68156
rect 113140 68184 113146 68196
rect 146478 68184 146484 68196
rect 113140 68156 146484 68184
rect 113140 68144 113146 68156
rect 146478 68144 146484 68156
rect 146536 68144 146542 68196
rect 162302 68144 162308 68196
rect 162360 68184 162366 68196
rect 182910 68184 182916 68196
rect 162360 68156 182916 68184
rect 162360 68144 162366 68156
rect 182910 68144 182916 68156
rect 182968 68144 182974 68196
rect 103054 68076 103060 68128
rect 103112 68116 103118 68128
rect 138382 68116 138388 68128
rect 103112 68088 138388 68116
rect 103112 68076 103118 68088
rect 138382 68076 138388 68088
rect 138440 68076 138446 68128
rect 160370 68076 160376 68128
rect 160428 68116 160434 68128
rect 161382 68116 161388 68128
rect 160428 68088 161388 68116
rect 160428 68076 160434 68088
rect 161382 68076 161388 68088
rect 161440 68076 161446 68128
rect 168098 68076 168104 68128
rect 168156 68116 168162 68128
rect 202046 68116 202052 68128
rect 168156 68088 202052 68116
rect 168156 68076 168162 68088
rect 202046 68076 202052 68088
rect 202104 68076 202110 68128
rect 107562 68008 107568 68060
rect 107620 68048 107626 68060
rect 135530 68048 135536 68060
rect 107620 68020 135536 68048
rect 107620 68008 107626 68020
rect 135530 68008 135536 68020
rect 135588 68008 135594 68060
rect 158438 68008 158444 68060
rect 158496 68048 158502 68060
rect 160462 68048 160468 68060
rect 158496 68020 160468 68048
rect 158496 68008 158502 68020
rect 160462 68008 160468 68020
rect 160520 68008 160526 68060
rect 162762 68008 162768 68060
rect 162820 68048 162826 68060
rect 171962 68048 171968 68060
rect 162820 68020 171968 68048
rect 162820 68008 162826 68020
rect 171962 68008 171968 68020
rect 172020 68008 172026 68060
rect 161842 67940 161848 67992
rect 161900 67980 161906 67992
rect 171870 67980 171876 67992
rect 161900 67952 171876 67980
rect 161900 67940 161906 67952
rect 171870 67940 171876 67952
rect 171928 67940 171934 67992
rect 160554 67872 160560 67924
rect 160612 67912 160618 67924
rect 161290 67912 161296 67924
rect 160612 67884 161296 67912
rect 160612 67872 160618 67884
rect 161290 67872 161296 67884
rect 161348 67872 161354 67924
rect 159082 67600 159088 67652
rect 159140 67640 159146 67652
rect 160002 67640 160008 67652
rect 159140 67612 160008 67640
rect 159140 67600 159146 67612
rect 160002 67600 160008 67612
rect 160060 67600 160066 67652
rect 167362 67600 167368 67652
rect 167420 67640 167426 67652
rect 168098 67640 168104 67652
rect 167420 67612 168104 67640
rect 167420 67600 167426 67612
rect 168098 67600 168104 67612
rect 168156 67600 168162 67652
rect 96430 67532 96436 67584
rect 96488 67572 96494 67584
rect 141050 67572 141056 67584
rect 96488 67544 141056 67572
rect 96488 67532 96494 67544
rect 141050 67532 141056 67544
rect 141108 67532 141114 67584
rect 168190 67532 168196 67584
rect 168248 67572 168254 67584
rect 217502 67572 217508 67584
rect 168248 67544 217508 67572
rect 168248 67532 168254 67544
rect 217502 67532 217508 67544
rect 217560 67572 217566 67584
rect 580626 67572 580632 67584
rect 217560 67544 580632 67572
rect 217560 67532 217566 67544
rect 580626 67532 580632 67544
rect 580684 67532 580690 67584
rect 109954 67464 109960 67516
rect 110012 67504 110018 67516
rect 143994 67504 144000 67516
rect 110012 67476 144000 67504
rect 110012 67464 110018 67476
rect 143994 67464 144000 67476
rect 144052 67464 144058 67516
rect 176654 67464 176660 67516
rect 176712 67504 176718 67516
rect 211614 67504 211620 67516
rect 176712 67476 211620 67504
rect 176712 67464 176718 67476
rect 211614 67464 211620 67476
rect 211672 67504 211678 67516
rect 212442 67504 212448 67516
rect 211672 67476 212448 67504
rect 211672 67464 211678 67476
rect 212442 67464 212448 67476
rect 212500 67464 212506 67516
rect 110046 67396 110052 67448
rect 110104 67436 110110 67448
rect 144270 67436 144276 67448
rect 110104 67408 144276 67436
rect 110104 67396 110110 67408
rect 144270 67396 144276 67408
rect 144328 67396 144334 67448
rect 163222 67396 163228 67448
rect 163280 67436 163286 67448
rect 198090 67436 198096 67448
rect 163280 67408 198096 67436
rect 163280 67396 163286 67408
rect 198090 67396 198096 67408
rect 198148 67396 198154 67448
rect 104618 67328 104624 67380
rect 104676 67368 104682 67380
rect 104676 67340 135392 67368
rect 104676 67328 104682 67340
rect 104710 67260 104716 67312
rect 104768 67300 104774 67312
rect 135254 67300 135260 67312
rect 104768 67272 135260 67300
rect 104768 67260 104774 67272
rect 135254 67260 135260 67272
rect 135312 67260 135318 67312
rect 135364 67300 135392 67340
rect 135438 67328 135444 67380
rect 135496 67368 135502 67380
rect 136082 67368 136088 67380
rect 135496 67340 136088 67368
rect 135496 67328 135502 67340
rect 136082 67328 136088 67340
rect 136140 67328 136146 67380
rect 137002 67328 137008 67380
rect 137060 67368 137066 67380
rect 137278 67368 137284 67380
rect 137060 67340 137284 67368
rect 137060 67328 137066 67340
rect 137278 67328 137284 67340
rect 137336 67328 137342 67380
rect 138658 67328 138664 67380
rect 138716 67368 138722 67380
rect 139302 67368 139308 67380
rect 138716 67340 139308 67368
rect 138716 67328 138722 67340
rect 139302 67328 139308 67340
rect 139360 67328 139366 67380
rect 139394 67328 139400 67380
rect 139452 67368 139458 67380
rect 140498 67368 140504 67380
rect 139452 67340 140504 67368
rect 139452 67328 139458 67340
rect 140498 67328 140504 67340
rect 140556 67328 140562 67380
rect 174078 67328 174084 67380
rect 174136 67368 174142 67380
rect 208670 67368 208676 67380
rect 174136 67340 208676 67368
rect 174136 67328 174142 67340
rect 208670 67328 208676 67340
rect 208728 67328 208734 67380
rect 138014 67300 138020 67312
rect 135364 67272 138020 67300
rect 138014 67260 138020 67272
rect 138072 67260 138078 67312
rect 160278 67260 160284 67312
rect 160336 67300 160342 67312
rect 194778 67300 194784 67312
rect 160336 67272 194784 67300
rect 160336 67260 160342 67272
rect 194778 67260 194784 67272
rect 194836 67260 194842 67312
rect 108942 67192 108948 67244
rect 109000 67232 109006 67244
rect 142338 67232 142344 67244
rect 109000 67204 142344 67232
rect 109000 67192 109006 67204
rect 142338 67192 142344 67204
rect 142396 67232 142402 67244
rect 142798 67232 142804 67244
rect 142396 67204 142804 67232
rect 142396 67192 142402 67204
rect 142798 67192 142804 67204
rect 142856 67192 142862 67244
rect 164510 67192 164516 67244
rect 164568 67232 164574 67244
rect 199010 67232 199016 67244
rect 164568 67204 199016 67232
rect 164568 67192 164574 67204
rect 199010 67192 199016 67204
rect 199068 67192 199074 67244
rect 110414 67124 110420 67176
rect 110472 67164 110478 67176
rect 112530 67164 112536 67176
rect 110472 67136 112536 67164
rect 110472 67124 110478 67136
rect 112530 67124 112536 67136
rect 112588 67164 112594 67176
rect 147122 67164 147128 67176
rect 112588 67136 147128 67164
rect 112588 67124 112594 67136
rect 147122 67124 147128 67136
rect 147180 67124 147186 67176
rect 164602 67124 164608 67176
rect 164660 67164 164666 67176
rect 199102 67164 199108 67176
rect 164660 67136 199108 67164
rect 164660 67124 164666 67136
rect 199102 67124 199108 67136
rect 199160 67124 199166 67176
rect 137186 67096 137192 67108
rect 103486 67068 137192 67096
rect 26234 66852 26240 66904
rect 26292 66892 26298 66904
rect 103146 66892 103152 66904
rect 26292 66864 103152 66892
rect 26292 66852 26298 66864
rect 103146 66852 103152 66864
rect 103204 66892 103210 66904
rect 103486 66892 103514 67068
rect 137186 67056 137192 67068
rect 137244 67056 137250 67108
rect 138014 67056 138020 67108
rect 138072 67096 138078 67108
rect 138750 67096 138756 67108
rect 138072 67068 138756 67096
rect 138072 67056 138078 67068
rect 138750 67056 138756 67068
rect 138808 67056 138814 67108
rect 163682 67056 163688 67108
rect 163740 67096 163746 67108
rect 164142 67096 164148 67108
rect 163740 67068 164148 67096
rect 163740 67056 163746 67068
rect 164142 67056 164148 67068
rect 164200 67096 164206 67108
rect 197722 67096 197728 67108
rect 164200 67068 197728 67096
rect 164200 67056 164206 67068
rect 197722 67056 197728 67068
rect 197780 67056 197786 67108
rect 104342 66988 104348 67040
rect 104400 67028 104406 67040
rect 137278 67028 137284 67040
rect 104400 67000 137284 67028
rect 104400 66988 104406 67000
rect 137278 66988 137284 67000
rect 137336 66988 137342 67040
rect 170398 66988 170404 67040
rect 170456 67028 170462 67040
rect 204530 67028 204536 67040
rect 170456 67000 204536 67028
rect 170456 66988 170462 67000
rect 204530 66988 204536 67000
rect 204588 66988 204594 67040
rect 107378 66920 107384 66972
rect 107436 66960 107442 66972
rect 135162 66960 135168 66972
rect 107436 66932 135168 66960
rect 107436 66920 107442 66932
rect 135162 66920 135168 66932
rect 135220 66920 135226 66972
rect 135254 66920 135260 66972
rect 135312 66960 135318 66972
rect 138658 66960 138664 66972
rect 135312 66932 138664 66960
rect 135312 66920 135318 66932
rect 138658 66920 138664 66932
rect 138716 66920 138722 66972
rect 166902 66920 166908 66972
rect 166960 66960 166966 66972
rect 200206 66960 200212 66972
rect 166960 66932 200212 66960
rect 166960 66920 166966 66932
rect 200206 66920 200212 66932
rect 200264 66920 200270 66972
rect 212442 66920 212448 66972
rect 212500 66960 212506 66972
rect 235994 66960 236000 66972
rect 212500 66932 236000 66960
rect 212500 66920 212506 66932
rect 235994 66920 236000 66932
rect 236052 66920 236058 66972
rect 103204 66864 103514 66892
rect 103204 66852 103210 66864
rect 116486 66852 116492 66904
rect 116544 66892 116550 66904
rect 148134 66892 148140 66904
rect 116544 66864 148140 66892
rect 116544 66852 116550 66864
rect 148134 66852 148140 66864
rect 148192 66892 148198 66904
rect 148318 66892 148324 66904
rect 148192 66864 148324 66892
rect 148192 66852 148198 66864
rect 148318 66852 148324 66864
rect 148376 66852 148382 66904
rect 150158 66852 150164 66904
rect 150216 66892 150222 66904
rect 503714 66892 503720 66904
rect 150216 66864 503720 66892
rect 150216 66852 150222 66864
rect 503714 66852 503720 66864
rect 503772 66852 503778 66904
rect 103422 66784 103428 66836
rect 103480 66824 103486 66836
rect 134334 66824 134340 66836
rect 103480 66796 134340 66824
rect 103480 66784 103486 66796
rect 134334 66784 134340 66796
rect 134392 66784 134398 66836
rect 108758 66716 108764 66768
rect 108816 66756 108822 66768
rect 139394 66756 139400 66768
rect 108816 66728 139400 66756
rect 108816 66716 108822 66728
rect 139394 66716 139400 66728
rect 139452 66716 139458 66768
rect 106090 66648 106096 66700
rect 106148 66688 106154 66700
rect 135438 66688 135444 66700
rect 106148 66660 135444 66688
rect 106148 66648 106154 66660
rect 135438 66648 135444 66660
rect 135496 66648 135502 66700
rect 135162 66580 135168 66632
rect 135220 66620 135226 66632
rect 140682 66620 140688 66632
rect 135220 66592 140688 66620
rect 135220 66580 135226 66592
rect 140682 66580 140688 66592
rect 140740 66580 140746 66632
rect 170398 66308 170404 66360
rect 170456 66348 170462 66360
rect 170950 66348 170956 66360
rect 170456 66320 170956 66348
rect 170456 66308 170462 66320
rect 170950 66308 170956 66320
rect 171008 66308 171014 66360
rect 346394 66280 346400 66292
rect 142126 66252 346400 66280
rect 120810 66172 120816 66224
rect 120868 66212 120874 66224
rect 141142 66212 141148 66224
rect 120868 66184 141148 66212
rect 120868 66172 120874 66184
rect 141142 66172 141148 66184
rect 141200 66212 141206 66224
rect 142126 66212 142154 66252
rect 346394 66240 346400 66252
rect 346452 66240 346458 66292
rect 141200 66184 142154 66212
rect 141200 66172 141206 66184
rect 142614 66172 142620 66224
rect 142672 66212 142678 66224
rect 142890 66212 142896 66224
rect 142672 66184 142896 66212
rect 142672 66172 142678 66184
rect 142890 66172 142896 66184
rect 142948 66172 142954 66224
rect 158898 66172 158904 66224
rect 158956 66212 158962 66224
rect 219802 66212 219808 66224
rect 158956 66184 219808 66212
rect 158956 66172 158962 66184
rect 219802 66172 219808 66184
rect 219860 66172 219866 66224
rect 102778 66104 102784 66156
rect 102836 66144 102842 66156
rect 142706 66144 142712 66156
rect 102836 66116 142712 66144
rect 102836 66104 102842 66116
rect 142706 66104 142712 66116
rect 142764 66144 142770 66156
rect 143442 66144 143448 66156
rect 142764 66116 143448 66144
rect 142764 66104 142770 66116
rect 143442 66104 143448 66116
rect 143500 66104 143506 66156
rect 156322 66104 156328 66156
rect 156380 66144 156386 66156
rect 216674 66144 216680 66156
rect 156380 66116 216680 66144
rect 156380 66104 156386 66116
rect 216674 66104 216680 66116
rect 216732 66104 216738 66156
rect 116210 66036 116216 66088
rect 116268 66076 116274 66088
rect 155586 66076 155592 66088
rect 116268 66048 155592 66076
rect 116268 66036 116274 66048
rect 155586 66036 155592 66048
rect 155644 66036 155650 66088
rect 170030 66036 170036 66088
rect 170088 66076 170094 66088
rect 209774 66076 209780 66088
rect 170088 66048 209780 66076
rect 170088 66036 170094 66048
rect 209774 66036 209780 66048
rect 209832 66036 209838 66088
rect 117222 65968 117228 66020
rect 117280 66008 117286 66020
rect 153378 66008 153384 66020
rect 117280 65980 153384 66008
rect 117280 65968 117286 65980
rect 153378 65968 153384 65980
rect 153436 65968 153442 66020
rect 164418 65968 164424 66020
rect 164476 66008 164482 66020
rect 203242 66008 203248 66020
rect 164476 65980 203248 66008
rect 164476 65968 164482 65980
rect 203242 65968 203248 65980
rect 203300 65968 203306 66020
rect 100018 65900 100024 65952
rect 100076 65940 100082 65952
rect 134886 65940 134892 65952
rect 100076 65912 134892 65940
rect 100076 65900 100082 65912
rect 134886 65900 134892 65912
rect 134944 65900 134950 65952
rect 158070 65900 158076 65952
rect 158128 65940 158134 65952
rect 192110 65940 192116 65952
rect 158128 65912 192116 65940
rect 158128 65900 158134 65912
rect 192110 65900 192116 65912
rect 192168 65940 192174 65952
rect 193122 65940 193128 65952
rect 192168 65912 193128 65940
rect 192168 65900 192174 65912
rect 193122 65900 193128 65912
rect 193180 65900 193186 65952
rect 101306 65832 101312 65884
rect 101364 65872 101370 65884
rect 136450 65872 136456 65884
rect 101364 65844 136456 65872
rect 101364 65832 101370 65844
rect 136450 65832 136456 65844
rect 136508 65872 136514 65884
rect 146938 65872 146944 65884
rect 136508 65844 146944 65872
rect 136508 65832 136514 65844
rect 146938 65832 146944 65844
rect 146996 65832 147002 65884
rect 173802 65832 173808 65884
rect 173860 65872 173866 65884
rect 208394 65872 208400 65884
rect 173860 65844 208400 65872
rect 173860 65832 173866 65844
rect 208394 65832 208400 65844
rect 208452 65832 208458 65884
rect 99926 65764 99932 65816
rect 99984 65804 99990 65816
rect 133046 65804 133052 65816
rect 99984 65776 133052 65804
rect 99984 65764 99990 65776
rect 133046 65764 133052 65776
rect 133104 65764 133110 65816
rect 153930 65764 153936 65816
rect 153988 65804 153994 65816
rect 188338 65804 188344 65816
rect 153988 65776 188344 65804
rect 153988 65764 153994 65776
rect 188338 65764 188344 65776
rect 188396 65764 188402 65816
rect 105354 65696 105360 65748
rect 105412 65736 105418 65748
rect 138198 65736 138204 65748
rect 105412 65708 138204 65736
rect 105412 65696 105418 65708
rect 138198 65696 138204 65708
rect 138256 65696 138262 65748
rect 167178 65696 167184 65748
rect 167236 65736 167242 65748
rect 168282 65736 168288 65748
rect 167236 65708 168288 65736
rect 167236 65696 167242 65708
rect 168282 65696 168288 65708
rect 168340 65736 168346 65748
rect 200666 65736 200672 65748
rect 168340 65708 200672 65736
rect 168340 65696 168346 65708
rect 200666 65696 200672 65708
rect 200724 65696 200730 65748
rect 102042 65628 102048 65680
rect 102100 65668 102106 65680
rect 134150 65668 134156 65680
rect 102100 65640 134156 65668
rect 102100 65628 102106 65640
rect 134150 65628 134156 65640
rect 134208 65628 134214 65680
rect 134886 65628 134892 65680
rect 134944 65668 134950 65680
rect 135898 65668 135904 65680
rect 134944 65640 135904 65668
rect 134944 65628 134950 65640
rect 135898 65628 135904 65640
rect 135956 65628 135962 65680
rect 161750 65628 161756 65680
rect 161808 65668 161814 65680
rect 189442 65668 189448 65680
rect 161808 65640 189448 65668
rect 161808 65628 161814 65640
rect 189442 65628 189448 65640
rect 189500 65628 189506 65680
rect 193122 65628 193128 65680
rect 193180 65668 193186 65680
rect 216674 65668 216680 65680
rect 193180 65640 216680 65668
rect 193180 65628 193186 65640
rect 216674 65628 216680 65640
rect 216732 65628 216738 65680
rect 151262 65600 151268 65612
rect 122806 65572 151268 65600
rect 35158 65492 35164 65544
rect 35216 65532 35222 65544
rect 118418 65532 118424 65544
rect 35216 65504 118424 65532
rect 35216 65492 35222 65504
rect 118418 65492 118424 65504
rect 118476 65532 118482 65544
rect 122806 65532 122834 65572
rect 151262 65560 151268 65572
rect 151320 65560 151326 65612
rect 167270 65560 167276 65612
rect 167328 65600 167334 65612
rect 171134 65600 171140 65612
rect 167328 65572 171140 65600
rect 167328 65560 167334 65572
rect 171134 65560 171140 65572
rect 171192 65600 171198 65612
rect 201954 65600 201960 65612
rect 171192 65572 201960 65600
rect 171192 65560 171198 65572
rect 201954 65560 201960 65572
rect 202012 65560 202018 65612
rect 118476 65504 122834 65532
rect 118476 65492 118482 65504
rect 128446 65492 128452 65544
rect 128504 65532 128510 65544
rect 128998 65532 129004 65544
rect 128504 65504 129004 65532
rect 128504 65492 128510 65504
rect 128998 65492 129004 65504
rect 129056 65492 129062 65544
rect 143442 65492 143448 65544
rect 143500 65532 143506 65544
rect 438854 65532 438860 65544
rect 143500 65504 438860 65532
rect 143500 65492 143506 65504
rect 438854 65492 438860 65504
rect 438912 65492 438918 65544
rect 99834 65424 99840 65476
rect 99892 65464 99898 65476
rect 128464 65464 128492 65492
rect 139578 65464 139584 65476
rect 99892 65436 128492 65464
rect 132466 65436 139584 65464
rect 99892 65424 99898 65436
rect 132466 65408 132494 65436
rect 139578 65424 139584 65436
rect 139636 65424 139642 65476
rect 112162 65356 112168 65408
rect 112220 65396 112226 65408
rect 132466 65396 132500 65408
rect 112220 65368 132500 65396
rect 112220 65356 112226 65368
rect 132494 65356 132500 65368
rect 132552 65356 132558 65408
rect 134150 65356 134156 65408
rect 134208 65396 134214 65408
rect 134702 65396 134708 65408
rect 134208 65368 134708 65396
rect 134208 65356 134214 65368
rect 134702 65356 134708 65368
rect 134760 65356 134766 65408
rect 95142 65288 95148 65340
rect 95200 65328 95206 65340
rect 160186 65328 160192 65340
rect 95200 65300 160192 65328
rect 95200 65288 95206 65300
rect 160186 65288 160192 65300
rect 160244 65288 160250 65340
rect 121822 65220 121828 65272
rect 121880 65260 121886 65272
rect 142890 65260 142896 65272
rect 121880 65232 142896 65260
rect 121880 65220 121886 65232
rect 142890 65220 142896 65232
rect 142948 65220 142954 65272
rect 3142 64812 3148 64864
rect 3200 64852 3206 64864
rect 158438 64852 158444 64864
rect 3200 64824 158444 64852
rect 3200 64812 3206 64824
rect 158438 64812 158444 64824
rect 158496 64812 158502 64864
rect 169846 64812 169852 64864
rect 169904 64852 169910 64864
rect 171042 64852 171048 64864
rect 169904 64824 171048 64852
rect 169904 64812 169910 64824
rect 171042 64812 171048 64824
rect 171100 64812 171106 64864
rect 171226 64812 171232 64864
rect 171284 64852 171290 64864
rect 171870 64852 171876 64864
rect 171284 64824 171876 64852
rect 171284 64812 171290 64824
rect 171870 64812 171876 64824
rect 171928 64812 171934 64864
rect 175458 64812 175464 64864
rect 175516 64852 175522 64864
rect 175918 64852 175924 64864
rect 175516 64824 175924 64852
rect 175516 64812 175522 64824
rect 175918 64812 175924 64824
rect 175976 64852 175982 64864
rect 212534 64852 212540 64864
rect 175976 64824 212540 64852
rect 175976 64812 175982 64824
rect 212534 64812 212540 64824
rect 212592 64812 212598 64864
rect 96338 64744 96344 64796
rect 96396 64784 96402 64796
rect 146662 64784 146668 64796
rect 96396 64756 146668 64784
rect 96396 64744 96402 64756
rect 146662 64744 146668 64756
rect 146720 64744 146726 64796
rect 169938 64744 169944 64796
rect 169996 64784 170002 64796
rect 205726 64784 205732 64796
rect 169996 64756 205732 64784
rect 169996 64744 170002 64756
rect 205726 64744 205732 64756
rect 205784 64744 205790 64796
rect 118602 64676 118608 64728
rect 118660 64716 118666 64728
rect 153746 64716 153752 64728
rect 118660 64688 153752 64716
rect 118660 64676 118666 64688
rect 153746 64676 153752 64688
rect 153804 64676 153810 64728
rect 165798 64676 165804 64728
rect 165856 64716 165862 64728
rect 200850 64716 200856 64728
rect 165856 64688 200856 64716
rect 165856 64676 165862 64688
rect 200850 64676 200856 64688
rect 200908 64676 200914 64728
rect 100570 64608 100576 64660
rect 100628 64648 100634 64660
rect 134610 64648 134616 64660
rect 100628 64620 134616 64648
rect 100628 64608 100634 64620
rect 134610 64608 134616 64620
rect 134668 64608 134674 64660
rect 173986 64608 173992 64660
rect 174044 64648 174050 64660
rect 175182 64648 175188 64660
rect 174044 64620 175188 64648
rect 174044 64608 174050 64620
rect 175182 64608 175188 64620
rect 175240 64648 175246 64660
rect 208762 64648 208768 64660
rect 175240 64620 208768 64648
rect 175240 64608 175246 64620
rect 208762 64608 208768 64620
rect 208820 64608 208826 64660
rect 106182 64540 106188 64592
rect 106240 64580 106246 64592
rect 140038 64580 140044 64592
rect 106240 64552 140044 64580
rect 106240 64540 106246 64552
rect 140038 64540 140044 64552
rect 140096 64540 140102 64592
rect 171870 64540 171876 64592
rect 171928 64580 171934 64592
rect 205910 64580 205916 64592
rect 171928 64552 205916 64580
rect 171928 64540 171934 64552
rect 205910 64540 205916 64552
rect 205968 64540 205974 64592
rect 100662 64472 100668 64524
rect 100720 64512 100726 64524
rect 132862 64512 132868 64524
rect 100720 64484 132868 64512
rect 100720 64472 100726 64484
rect 132862 64472 132868 64484
rect 132920 64512 132926 64524
rect 133782 64512 133788 64524
rect 132920 64484 133788 64512
rect 132920 64472 132926 64484
rect 133782 64472 133788 64484
rect 133840 64472 133846 64524
rect 173250 64472 173256 64524
rect 173308 64512 173314 64524
rect 173802 64512 173808 64524
rect 173308 64484 173808 64512
rect 173308 64472 173314 64484
rect 173802 64472 173808 64484
rect 173860 64512 173866 64524
rect 207014 64512 207020 64524
rect 173860 64484 207020 64512
rect 173860 64472 173866 64484
rect 207014 64472 207020 64484
rect 207072 64472 207078 64524
rect 104250 64404 104256 64456
rect 104308 64444 104314 64456
rect 136818 64444 136824 64456
rect 104308 64416 136824 64444
rect 104308 64404 104314 64416
rect 136818 64404 136824 64416
rect 136876 64404 136882 64456
rect 161658 64404 161664 64456
rect 161716 64444 161722 64456
rect 196066 64444 196072 64456
rect 161716 64416 196072 64444
rect 161716 64404 161722 64416
rect 196066 64404 196072 64416
rect 196124 64404 196130 64456
rect 122098 64336 122104 64388
rect 122156 64376 122162 64388
rect 154114 64376 154120 64388
rect 122156 64348 154120 64376
rect 122156 64336 122162 64348
rect 154114 64336 154120 64348
rect 154172 64336 154178 64388
rect 171042 64336 171048 64388
rect 171100 64376 171106 64388
rect 203886 64376 203892 64388
rect 171100 64348 203892 64376
rect 171100 64336 171106 64348
rect 203886 64336 203892 64348
rect 203944 64336 203950 64388
rect 128354 64268 128360 64320
rect 128412 64308 128418 64320
rect 207566 64308 207572 64320
rect 128412 64280 207572 64308
rect 128412 64268 128418 64280
rect 207566 64268 207572 64280
rect 207624 64268 207630 64320
rect 105998 64200 106004 64252
rect 106056 64240 106062 64252
rect 137830 64240 137836 64252
rect 106056 64212 137836 64240
rect 106056 64200 106062 64212
rect 137830 64200 137836 64212
rect 137888 64200 137894 64252
rect 143994 64200 144000 64252
rect 144052 64240 144058 64252
rect 278774 64240 278780 64252
rect 144052 64212 278780 64240
rect 144052 64200 144058 64212
rect 278774 64200 278780 64212
rect 278832 64200 278838 64252
rect 136818 64132 136824 64184
rect 136876 64172 136882 64184
rect 144914 64172 144920 64184
rect 136876 64144 144920 64172
rect 136876 64132 136882 64144
rect 144914 64132 144920 64144
rect 144972 64132 144978 64184
rect 154850 64132 154856 64184
rect 154908 64172 154914 64184
rect 154908 64144 157334 64172
rect 154908 64132 154914 64144
rect 157306 64036 157334 64144
rect 189074 64132 189080 64184
rect 189132 64172 189138 64184
rect 488534 64172 488540 64184
rect 189132 64144 488540 64172
rect 189132 64132 189138 64144
rect 488534 64132 488540 64144
rect 488592 64132 488598 64184
rect 162854 64064 162860 64116
rect 162912 64104 162918 64116
rect 163038 64104 163044 64116
rect 162912 64076 163044 64104
rect 162912 64064 162918 64076
rect 163038 64064 163044 64076
rect 163096 64104 163102 64116
rect 191282 64104 191288 64116
rect 163096 64076 191288 64104
rect 163096 64064 163102 64076
rect 191282 64064 191288 64076
rect 191340 64064 191346 64116
rect 165430 64036 165436 64048
rect 157306 64008 165436 64036
rect 165430 63996 165436 64008
rect 165488 64036 165494 64048
rect 189258 64036 189264 64048
rect 165488 64008 189264 64036
rect 165488 63996 165494 64008
rect 189258 63996 189264 64008
rect 189316 63996 189322 64048
rect 157702 63928 157708 63980
rect 157760 63968 157766 63980
rect 189074 63968 189080 63980
rect 157760 63940 189080 63968
rect 157760 63928 157766 63940
rect 189074 63928 189080 63940
rect 189132 63928 189138 63980
rect 96154 63452 96160 63504
rect 96212 63492 96218 63504
rect 143074 63492 143080 63504
rect 96212 63464 143080 63492
rect 96212 63452 96218 63464
rect 143074 63452 143080 63464
rect 143132 63452 143138 63504
rect 154022 63452 154028 63504
rect 154080 63492 154086 63504
rect 580350 63492 580356 63504
rect 154080 63464 580356 63492
rect 154080 63452 154086 63464
rect 580350 63452 580356 63464
rect 580408 63452 580414 63504
rect 97166 63384 97172 63436
rect 97224 63424 97230 63436
rect 139118 63424 139124 63436
rect 97224 63396 139124 63424
rect 97224 63384 97230 63396
rect 139118 63384 139124 63396
rect 139176 63384 139182 63436
rect 156874 63384 156880 63436
rect 156932 63424 156938 63436
rect 580534 63424 580540 63436
rect 156932 63396 580540 63424
rect 156932 63384 156938 63396
rect 580534 63384 580540 63396
rect 580592 63384 580598 63436
rect 100478 63316 100484 63368
rect 100536 63356 100542 63368
rect 141418 63356 141424 63368
rect 100536 63328 141424 63356
rect 100536 63316 100542 63328
rect 141418 63316 141424 63328
rect 141476 63316 141482 63368
rect 156230 63316 156236 63368
rect 156288 63356 156294 63368
rect 215662 63356 215668 63368
rect 156288 63328 215668 63356
rect 156288 63316 156294 63328
rect 215662 63316 215668 63328
rect 215720 63316 215726 63368
rect 96522 63248 96528 63300
rect 96580 63288 96586 63300
rect 134242 63288 134248 63300
rect 96580 63260 134248 63288
rect 96580 63248 96586 63260
rect 134242 63248 134248 63260
rect 134300 63248 134306 63300
rect 161474 63248 161480 63300
rect 161532 63288 161538 63300
rect 219526 63288 219532 63300
rect 161532 63260 219532 63288
rect 161532 63248 161538 63260
rect 219526 63248 219532 63260
rect 219584 63248 219590 63300
rect 162486 63180 162492 63232
rect 162544 63220 162550 63232
rect 210050 63220 210056 63232
rect 162544 63192 210056 63220
rect 162544 63180 162550 63192
rect 210050 63180 210056 63192
rect 210108 63180 210114 63232
rect 167914 63112 167920 63164
rect 167972 63152 167978 63164
rect 210510 63152 210516 63164
rect 167972 63124 210516 63152
rect 167972 63112 167978 63124
rect 210510 63112 210516 63124
rect 210568 63112 210574 63164
rect 164326 63044 164332 63096
rect 164384 63084 164390 63096
rect 165522 63084 165528 63096
rect 164384 63056 165528 63084
rect 164384 63044 164390 63056
rect 165522 63044 165528 63056
rect 165580 63084 165586 63096
rect 206278 63084 206284 63096
rect 165580 63056 206284 63084
rect 165580 63044 165586 63056
rect 206278 63044 206284 63056
rect 206336 63044 206342 63096
rect 167086 62976 167092 63028
rect 167144 63016 167150 63028
rect 208854 63016 208860 63028
rect 167144 62988 208860 63016
rect 167144 62976 167150 62988
rect 208854 62976 208860 62988
rect 208912 62976 208918 63028
rect 165706 62908 165712 62960
rect 165764 62948 165770 62960
rect 166902 62948 166908 62960
rect 165764 62920 166908 62948
rect 165764 62908 165770 62920
rect 166902 62908 166908 62920
rect 166960 62948 166966 62960
rect 207198 62948 207204 62960
rect 166960 62920 207204 62948
rect 166960 62908 166966 62920
rect 207198 62908 207204 62920
rect 207256 62908 207262 62960
rect 31018 62840 31024 62892
rect 31076 62880 31082 62892
rect 162854 62880 162860 62892
rect 31076 62852 162860 62880
rect 31076 62840 31082 62852
rect 162854 62840 162860 62852
rect 162912 62840 162918 62892
rect 168558 62840 168564 62892
rect 168616 62880 168622 62892
rect 182174 62880 182180 62892
rect 168616 62852 182180 62880
rect 168616 62840 168622 62852
rect 182174 62840 182180 62852
rect 182232 62880 182238 62892
rect 219434 62880 219440 62892
rect 182232 62852 219440 62880
rect 182232 62840 182238 62852
rect 219434 62840 219440 62852
rect 219492 62840 219498 62892
rect 142982 62772 142988 62824
rect 143040 62812 143046 62824
rect 430574 62812 430580 62824
rect 143040 62784 430580 62812
rect 143040 62772 143046 62784
rect 430574 62772 430580 62784
rect 430632 62772 430638 62824
rect 167730 62704 167736 62756
rect 167788 62744 167794 62756
rect 202230 62744 202236 62756
rect 167788 62716 202236 62744
rect 167788 62704 167794 62716
rect 202230 62704 202236 62716
rect 202288 62704 202294 62756
rect 134242 62092 134248 62144
rect 134300 62132 134306 62144
rect 134794 62132 134800 62144
rect 134300 62104 134800 62132
rect 134300 62092 134306 62104
rect 134794 62092 134800 62104
rect 134852 62092 134858 62144
rect 138842 62092 138848 62144
rect 138900 62132 138906 62144
rect 139118 62132 139124 62144
rect 138900 62104 139124 62132
rect 138900 62092 138906 62104
rect 139118 62092 139124 62104
rect 139176 62092 139182 62144
rect 158714 62024 158720 62076
rect 158772 62064 158778 62076
rect 193214 62064 193220 62076
rect 158772 62036 193220 62064
rect 158772 62024 158778 62036
rect 193214 62024 193220 62036
rect 193272 62064 193278 62076
rect 194502 62064 194508 62076
rect 193272 62036 194508 62064
rect 193272 62024 193278 62036
rect 194502 62024 194508 62036
rect 194560 62024 194566 62076
rect 155862 61956 155868 62008
rect 155920 61996 155926 62008
rect 186314 61996 186320 62008
rect 155920 61968 186320 61996
rect 155920 61956 155926 61968
rect 186314 61956 186320 61968
rect 186372 61956 186378 62008
rect 161198 61888 161204 61940
rect 161256 61928 161262 61940
rect 190546 61928 190552 61940
rect 161256 61900 190552 61928
rect 161256 61888 161262 61900
rect 190546 61888 190552 61900
rect 190604 61888 190610 61940
rect 137830 61412 137836 61464
rect 137888 61452 137894 61464
rect 385034 61452 385040 61464
rect 137888 61424 385040 61452
rect 137888 61412 137894 61424
rect 385034 61412 385040 61424
rect 385092 61412 385098 61464
rect 22738 61344 22744 61396
rect 22796 61384 22802 61396
rect 174814 61384 174820 61396
rect 22796 61356 174820 61384
rect 22796 61344 22802 61356
rect 174814 61344 174820 61356
rect 174872 61344 174878 61396
rect 194502 61344 194508 61396
rect 194560 61384 194566 61396
rect 558178 61384 558184 61396
rect 194560 61356 558184 61384
rect 194560 61344 194566 61356
rect 558178 61344 558184 61356
rect 558236 61344 558242 61396
rect 160094 61208 160100 61260
rect 160152 61248 160158 61260
rect 161198 61248 161204 61260
rect 160152 61220 161204 61248
rect 160152 61208 160158 61220
rect 161198 61208 161204 61220
rect 161256 61208 161262 61260
rect 96062 60664 96068 60716
rect 96120 60704 96126 60716
rect 139946 60704 139952 60716
rect 96120 60676 139952 60704
rect 96120 60664 96126 60676
rect 139946 60664 139952 60676
rect 140004 60664 140010 60716
rect 168466 60664 168472 60716
rect 168524 60704 168530 60716
rect 219710 60704 219716 60716
rect 168524 60676 219716 60704
rect 168524 60664 168530 60676
rect 219710 60664 219716 60676
rect 219768 60704 219774 60716
rect 220722 60704 220728 60716
rect 219768 60676 220728 60704
rect 219768 60664 219774 60676
rect 220722 60664 220728 60676
rect 220780 60664 220786 60716
rect 93118 60052 93124 60104
rect 93176 60092 93182 60104
rect 167086 60092 167092 60104
rect 93176 60064 167092 60092
rect 93176 60052 93182 60064
rect 167086 60052 167092 60064
rect 167144 60052 167150 60104
rect 220722 60052 220728 60104
rect 220780 60092 220786 60104
rect 404354 60092 404360 60104
rect 220780 60064 404360 60092
rect 220780 60052 220786 60064
rect 404354 60052 404360 60064
rect 404412 60052 404418 60104
rect 48314 59984 48320 60036
rect 48372 60024 48378 60036
rect 96062 60024 96068 60036
rect 48372 59996 96068 60024
rect 48372 59984 48378 59996
rect 96062 59984 96068 59996
rect 96120 59984 96126 60036
rect 144454 59984 144460 60036
rect 144512 60024 144518 60036
rect 342254 60024 342260 60036
rect 144512 59996 342260 60024
rect 144512 59984 144518 59996
rect 342254 59984 342260 59996
rect 342312 59984 342318 60036
rect 169662 59304 169668 59356
rect 169720 59344 169726 59356
rect 203518 59344 203524 59356
rect 169720 59316 203524 59344
rect 169720 59304 169726 59316
rect 203518 59304 203524 59316
rect 203576 59344 203582 59356
rect 204162 59344 204168 59356
rect 203576 59316 204168 59344
rect 203576 59304 203582 59316
rect 204162 59304 204168 59316
rect 204220 59304 204226 59356
rect 166166 59236 166172 59288
rect 166224 59276 166230 59288
rect 201126 59276 201132 59288
rect 166224 59248 201132 59276
rect 166224 59236 166230 59248
rect 201126 59236 201132 59248
rect 201184 59276 201190 59288
rect 201402 59276 201408 59288
rect 201184 59248 201408 59276
rect 201184 59236 201190 59248
rect 201402 59236 201408 59248
rect 201460 59236 201466 59288
rect 201402 58692 201408 58744
rect 201460 58732 201466 58744
rect 251174 58732 251180 58744
rect 201460 58704 251180 58732
rect 201460 58692 201466 58704
rect 251174 58692 251180 58704
rect 251232 58692 251238 58744
rect 95234 58624 95240 58676
rect 95292 58664 95298 58676
rect 166258 58664 166264 58676
rect 95292 58636 166264 58664
rect 95292 58624 95298 58636
rect 166258 58624 166264 58636
rect 166316 58624 166322 58676
rect 204162 58624 204168 58676
rect 204220 58664 204226 58676
rect 510614 58664 510620 58676
rect 204220 58636 510620 58664
rect 204220 58624 204226 58636
rect 510614 58624 510620 58636
rect 510672 58624 510678 58676
rect 169754 57876 169760 57928
rect 169812 57916 169818 57928
rect 204898 57916 204904 57928
rect 169812 57888 204904 57916
rect 169812 57876 169818 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 155494 57808 155500 57860
rect 155552 57848 155558 57860
rect 189074 57848 189080 57860
rect 155552 57820 189080 57848
rect 155552 57808 155558 57820
rect 189074 57808 189080 57820
rect 189132 57848 189138 57860
rect 189534 57848 189540 57860
rect 189132 57820 189540 57848
rect 189132 57808 189138 57820
rect 189534 57808 189540 57820
rect 189592 57808 189598 57860
rect 204898 57264 204904 57316
rect 204956 57304 204962 57316
rect 231854 57304 231860 57316
rect 204956 57276 231860 57304
rect 204956 57264 204962 57276
rect 231854 57264 231860 57276
rect 231912 57264 231918 57316
rect 6914 57196 6920 57248
rect 6972 57236 6978 57248
rect 160094 57236 160100 57248
rect 6972 57208 160100 57236
rect 6972 57196 6978 57208
rect 160094 57196 160100 57208
rect 160152 57196 160158 57248
rect 189074 57196 189080 57248
rect 189132 57236 189138 57248
rect 560294 57236 560300 57248
rect 189132 57208 560300 57236
rect 189132 57196 189138 57208
rect 560294 57196 560300 57208
rect 560352 57196 560358 57248
rect 3418 56516 3424 56568
rect 3476 56556 3482 56568
rect 97258 56556 97264 56568
rect 3476 56528 97264 56556
rect 3476 56516 3482 56528
rect 97258 56516 97264 56528
rect 97316 56516 97322 56568
rect 155402 56516 155408 56568
rect 155460 56556 155466 56568
rect 214558 56556 214564 56568
rect 155460 56528 214564 56556
rect 155460 56516 155466 56528
rect 214558 56516 214564 56528
rect 214616 56516 214622 56568
rect 17954 55904 17960 55956
rect 18012 55944 18018 55956
rect 176102 55944 176108 55956
rect 18012 55916 176108 55944
rect 18012 55904 18018 55916
rect 176102 55904 176108 55916
rect 176160 55904 176166 55956
rect 214558 55904 214564 55956
rect 214616 55944 214622 55956
rect 376754 55944 376760 55956
rect 214616 55916 376760 55944
rect 214616 55904 214622 55916
rect 376754 55904 376760 55916
rect 376812 55904 376818 55956
rect 133782 55836 133788 55888
rect 133840 55876 133846 55888
rect 538214 55876 538220 55888
rect 133840 55848 538220 55876
rect 133840 55836 133846 55848
rect 538214 55836 538220 55848
rect 538272 55836 538278 55888
rect 101398 55156 101404 55208
rect 101456 55196 101462 55208
rect 135714 55196 135720 55208
rect 101456 55168 135720 55196
rect 101456 55156 101462 55168
rect 135714 55156 135720 55168
rect 135772 55156 135778 55208
rect 162946 55156 162952 55208
rect 163004 55196 163010 55208
rect 198274 55196 198280 55208
rect 163004 55168 198280 55196
rect 163004 55156 163010 55168
rect 198274 55156 198280 55168
rect 198332 55156 198338 55208
rect 145650 54544 145656 54596
rect 145708 54584 145714 54596
rect 224954 54584 224960 54596
rect 145708 54556 224960 54584
rect 145708 54544 145714 54556
rect 224954 54544 224960 54556
rect 225012 54544 225018 54596
rect 13814 54476 13820 54528
rect 13872 54516 13878 54528
rect 101398 54516 101404 54528
rect 13872 54488 101404 54516
rect 13872 54476 13878 54488
rect 101398 54476 101404 54488
rect 101456 54476 101462 54528
rect 198274 54476 198280 54528
rect 198332 54516 198338 54528
rect 400214 54516 400220 54528
rect 198332 54488 400220 54516
rect 198332 54476 198338 54488
rect 400214 54476 400220 54488
rect 400272 54476 400278 54528
rect 105446 53728 105452 53780
rect 105504 53768 105510 53780
rect 138566 53768 138572 53780
rect 105504 53740 138572 53768
rect 105504 53728 105510 53740
rect 138566 53728 138572 53740
rect 138624 53728 138630 53780
rect 141418 53116 141424 53168
rect 141476 53156 141482 53168
rect 205634 53156 205640 53168
rect 141476 53128 205640 53156
rect 141476 53116 141482 53128
rect 205634 53116 205640 53128
rect 205692 53116 205698 53168
rect 3510 53048 3516 53100
rect 3568 53088 3574 53100
rect 105446 53088 105452 53100
rect 3568 53060 105452 53088
rect 3568 53048 3574 53060
rect 105446 53048 105452 53060
rect 105504 53048 105510 53100
rect 149882 53048 149888 53100
rect 149940 53088 149946 53100
rect 469214 53088 469220 53100
rect 149940 53060 469220 53088
rect 149940 53048 149946 53060
rect 469214 53048 469220 53060
rect 469272 53048 469278 53100
rect 3418 52368 3424 52420
rect 3476 52408 3482 52420
rect 110322 52408 110328 52420
rect 3476 52380 110328 52408
rect 3476 52368 3482 52380
rect 110322 52368 110328 52380
rect 110380 52408 110386 52420
rect 138934 52408 138940 52420
rect 110380 52380 138940 52408
rect 110380 52368 110386 52380
rect 138934 52368 138940 52380
rect 138992 52368 138998 52420
rect 164234 52368 164240 52420
rect 164292 52408 164298 52420
rect 219618 52408 219624 52420
rect 164292 52380 219624 52408
rect 164292 52368 164298 52380
rect 219618 52368 219624 52380
rect 219676 52408 219682 52420
rect 220722 52408 220728 52420
rect 219676 52380 220728 52408
rect 219676 52368 219682 52380
rect 220722 52368 220728 52380
rect 220780 52368 220786 52420
rect 149790 51756 149796 51808
rect 149848 51796 149854 51808
rect 309134 51796 309140 51808
rect 149848 51768 309140 51796
rect 149848 51756 149854 51768
rect 309134 51756 309140 51768
rect 309192 51756 309198 51808
rect 220722 51688 220728 51740
rect 220780 51728 220786 51740
rect 563698 51728 563704 51740
rect 220780 51700 563704 51728
rect 220780 51688 220786 51700
rect 563698 51688 563704 51700
rect 563756 51688 563762 51740
rect 164050 51008 164056 51060
rect 164108 51048 164114 51060
rect 197446 51048 197452 51060
rect 164108 51020 197452 51048
rect 164108 51008 164114 51020
rect 197446 51008 197452 51020
rect 197504 51008 197510 51060
rect 149698 50396 149704 50448
rect 149756 50436 149762 50448
rect 304994 50436 305000 50448
rect 149756 50408 305000 50436
rect 149756 50396 149762 50408
rect 304994 50396 305000 50408
rect 305052 50396 305058 50448
rect 197446 50328 197452 50380
rect 197504 50368 197510 50380
rect 542998 50368 543004 50380
rect 197504 50340 543004 50368
rect 197504 50328 197510 50340
rect 542998 50328 543004 50340
rect 543056 50328 543062 50380
rect 3234 49648 3240 49700
rect 3292 49688 3298 49700
rect 162118 49688 162124 49700
rect 3292 49660 162124 49688
rect 3292 49648 3298 49660
rect 162118 49648 162124 49660
rect 162176 49648 162182 49700
rect 183462 49648 183468 49700
rect 183520 49688 183526 49700
rect 580166 49688 580172 49700
rect 183520 49660 580172 49688
rect 183520 49648 183526 49660
rect 580166 49648 580172 49660
rect 580224 49648 580230 49700
rect 140130 48968 140136 49020
rect 140188 49008 140194 49020
rect 373994 49008 374000 49020
rect 140188 48980 374000 49008
rect 140188 48968 140194 48980
rect 373994 48968 374000 48980
rect 374052 48968 374058 49020
rect 156138 48220 156144 48272
rect 156196 48260 156202 48272
rect 190638 48260 190644 48272
rect 156196 48232 190644 48260
rect 156196 48220 156202 48232
rect 190638 48220 190644 48232
rect 190696 48260 190702 48272
rect 191742 48260 191748 48272
rect 190696 48232 191748 48260
rect 190696 48220 190702 48232
rect 191742 48220 191748 48232
rect 191800 48220 191806 48272
rect 191742 47608 191748 47660
rect 191800 47648 191806 47660
rect 369854 47648 369860 47660
rect 191800 47620 369860 47648
rect 191800 47608 191806 47620
rect 369854 47608 369860 47620
rect 369912 47608 369918 47660
rect 137278 47540 137284 47592
rect 137336 47580 137342 47592
rect 442258 47580 442264 47592
rect 137336 47552 442264 47580
rect 137336 47540 137342 47552
rect 442258 47540 442264 47552
rect 442316 47540 442322 47592
rect 156046 46860 156052 46912
rect 156104 46900 156110 46912
rect 215662 46900 215668 46912
rect 156104 46872 215668 46900
rect 156104 46860 156110 46872
rect 215662 46860 215668 46872
rect 215720 46900 215726 46912
rect 216030 46900 216036 46912
rect 215720 46872 216036 46900
rect 215720 46860 215726 46872
rect 216030 46860 216036 46872
rect 216088 46860 216094 46912
rect 215662 46248 215668 46300
rect 215720 46288 215726 46300
rect 396074 46288 396080 46300
rect 215720 46260 396080 46288
rect 215720 46248 215726 46260
rect 396074 46248 396080 46260
rect 396132 46248 396138 46300
rect 134794 46180 134800 46232
rect 134852 46220 134858 46232
rect 324314 46220 324320 46232
rect 134852 46192 324320 46220
rect 134852 46180 134858 46192
rect 324314 46180 324320 46192
rect 324372 46180 324378 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 22738 45540 22744 45552
rect 3568 45512 22744 45540
rect 3568 45500 3574 45512
rect 22738 45500 22744 45512
rect 22796 45500 22802 45552
rect 147030 45500 147036 45552
rect 147088 45540 147094 45552
rect 579982 45540 579988 45552
rect 147088 45512 579988 45540
rect 147088 45500 147094 45512
rect 579982 45500 579988 45512
rect 580040 45500 580046 45552
rect 144362 43460 144368 43512
rect 144420 43500 144426 43512
rect 354674 43500 354680 43512
rect 144420 43472 354680 43500
rect 144420 43460 144426 43472
rect 354674 43460 354680 43472
rect 354732 43460 354738 43512
rect 140038 43392 140044 43444
rect 140096 43432 140102 43444
rect 456794 43432 456800 43444
rect 140096 43404 456800 43432
rect 140096 43392 140102 43404
rect 456794 43392 456800 43404
rect 456852 43392 456858 43444
rect 134702 42100 134708 42152
rect 134760 42140 134766 42152
rect 242894 42140 242900 42152
rect 134760 42112 242900 42140
rect 134760 42100 134766 42112
rect 242894 42100 242900 42112
rect 242952 42100 242958 42152
rect 161290 42032 161296 42084
rect 161348 42072 161354 42084
rect 521654 42072 521660 42084
rect 161348 42044 521660 42072
rect 161348 42032 161354 42044
rect 521654 42032 521660 42044
rect 521712 42032 521718 42084
rect 3510 41352 3516 41404
rect 3568 41392 3574 41404
rect 122190 41392 122196 41404
rect 3568 41364 122196 41392
rect 3568 41352 3574 41364
rect 122190 41352 122196 41364
rect 122248 41352 122254 41404
rect 185578 41352 185584 41404
rect 185636 41392 185642 41404
rect 580166 41392 580172 41404
rect 185636 41364 580172 41392
rect 185636 41352 185642 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 148318 40672 148324 40724
rect 148376 40712 148382 40724
rect 193214 40712 193220 40724
rect 148376 40684 193220 40712
rect 148376 40672 148382 40684
rect 193214 40672 193220 40684
rect 193272 40672 193278 40724
rect 161382 39312 161388 39364
rect 161440 39352 161446 39364
rect 578878 39352 578884 39364
rect 161440 39324 578884 39352
rect 161440 39312 161446 39324
rect 578878 39312 578884 39324
rect 578936 39312 578942 39364
rect 164142 37952 164148 38004
rect 164200 37992 164206 38004
rect 331214 37992 331220 38004
rect 164200 37964 331220 37992
rect 164200 37952 164206 37964
rect 331214 37952 331220 37964
rect 331272 37952 331278 38004
rect 137094 37884 137100 37936
rect 137152 37924 137158 37936
rect 389174 37924 389180 37936
rect 137152 37896 389180 37924
rect 137152 37884 137158 37896
rect 389174 37884 389180 37896
rect 389232 37884 389238 37936
rect 3142 37204 3148 37256
rect 3200 37244 3206 37256
rect 128446 37244 128452 37256
rect 3200 37216 128452 37244
rect 3200 37204 3206 37216
rect 128446 37204 128452 37216
rect 128504 37204 128510 37256
rect 155954 37204 155960 37256
rect 156012 37244 156018 37256
rect 197354 37244 197360 37256
rect 156012 37216 197360 37244
rect 156012 37204 156018 37216
rect 197354 37204 197360 37216
rect 197412 37244 197418 37256
rect 580166 37244 580172 37256
rect 197412 37216 580172 37244
rect 197412 37204 197418 37216
rect 580166 37204 580172 37216
rect 580224 37204 580230 37256
rect 165338 35232 165344 35284
rect 165396 35272 165402 35284
rect 247034 35272 247040 35284
rect 165396 35244 247040 35272
rect 165396 35232 165402 35244
rect 247034 35232 247040 35244
rect 247092 35232 247098 35284
rect 153930 35164 153936 35216
rect 153988 35204 153994 35216
rect 499574 35204 499580 35216
rect 153988 35176 499580 35204
rect 153988 35164 153994 35176
rect 499574 35164 499580 35176
rect 499632 35164 499638 35216
rect 168190 33736 168196 33788
rect 168248 33776 168254 33788
rect 423674 33776 423680 33788
rect 168248 33748 423680 33776
rect 168248 33736 168254 33748
rect 423674 33736 423680 33748
rect 423732 33736 423738 33788
rect 158530 33056 158536 33108
rect 158588 33096 158594 33108
rect 580166 33096 580172 33108
rect 158588 33068 580172 33096
rect 158588 33056 158594 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3142 32988 3148 33040
rect 3200 33028 3206 33040
rect 177298 33028 177304 33040
rect 3200 33000 177304 33028
rect 3200 32988 3206 33000
rect 177298 32988 177304 33000
rect 177356 32988 177362 33040
rect 168282 31016 168288 31068
rect 168340 31056 168346 31068
rect 495434 31056 495440 31068
rect 168340 31028 495440 31056
rect 168340 31016 168346 31028
rect 495434 31016 495440 31028
rect 495492 31016 495498 31068
rect 162670 29656 162676 29708
rect 162728 29696 162734 29708
rect 357434 29696 357440 29708
rect 162728 29668 357440 29696
rect 162728 29656 162734 29668
rect 357434 29656 357440 29668
rect 357492 29656 357498 29708
rect 133138 29588 133144 29640
rect 133196 29628 133202 29640
rect 507854 29628 507860 29640
rect 133196 29600 507860 29628
rect 133196 29588 133202 29600
rect 507854 29588 507860 29600
rect 507912 29588 507918 29640
rect 3142 28908 3148 28960
rect 3200 28948 3206 28960
rect 147766 28948 147772 28960
rect 3200 28920 147772 28948
rect 3200 28908 3206 28920
rect 147766 28908 147772 28920
rect 147824 28908 147830 28960
rect 170950 28296 170956 28348
rect 171008 28336 171014 28348
rect 296714 28336 296720 28348
rect 171008 28308 296720 28336
rect 171008 28296 171014 28308
rect 296714 28296 296720 28308
rect 296772 28296 296778 28348
rect 144270 28228 144276 28280
rect 144328 28268 144334 28280
rect 571334 28268 571340 28280
rect 144328 28240 571340 28268
rect 144328 28228 144334 28240
rect 571334 28228 571340 28240
rect 571392 28228 571398 28280
rect 175182 26868 175188 26920
rect 175240 26908 175246 26920
rect 480254 26908 480260 26920
rect 175240 26880 480260 26908
rect 175240 26868 175246 26880
rect 480254 26868 480260 26880
rect 480312 26868 480318 26920
rect 166994 26256 167000 26308
rect 167052 26296 167058 26308
rect 171870 26296 171876 26308
rect 167052 26268 171876 26296
rect 167052 26256 167058 26268
rect 171870 26256 171876 26268
rect 171928 26256 171934 26308
rect 173802 25576 173808 25628
rect 173860 25616 173866 25628
rect 262214 25616 262220 25628
rect 173860 25588 262220 25616
rect 173860 25576 173866 25588
rect 262214 25576 262220 25588
rect 262272 25576 262278 25628
rect 155862 25508 155868 25560
rect 155920 25548 155926 25560
rect 575474 25548 575480 25560
rect 155920 25520 575480 25548
rect 155920 25508 155926 25520
rect 575474 25508 575480 25520
rect 575532 25508 575538 25560
rect 3050 24760 3056 24812
rect 3108 24800 3114 24812
rect 35158 24800 35164 24812
rect 3108 24772 35164 24800
rect 3108 24760 3114 24772
rect 35158 24760 35164 24772
rect 35216 24760 35222 24812
rect 184198 24760 184204 24812
rect 184256 24800 184262 24812
rect 580166 24800 580172 24812
rect 184256 24772 580172 24800
rect 184256 24760 184262 24772
rect 580166 24760 580172 24772
rect 580224 24760 580230 24812
rect 171042 22788 171048 22840
rect 171100 22828 171106 22840
rect 350534 22828 350540 22840
rect 171100 22800 350540 22828
rect 171100 22788 171106 22800
rect 350534 22788 350540 22800
rect 350592 22788 350598 22840
rect 138750 22720 138756 22772
rect 138808 22760 138814 22772
rect 392578 22760 392584 22772
rect 138808 22732 392584 22760
rect 138808 22720 138814 22732
rect 392578 22720 392584 22732
rect 392636 22720 392642 22772
rect 144178 21428 144184 21480
rect 144236 21468 144242 21480
rect 320174 21468 320180 21480
rect 144236 21440 320180 21468
rect 144236 21428 144242 21440
rect 320174 21428 320180 21440
rect 320232 21428 320238 21480
rect 138842 21360 138848 21412
rect 138900 21400 138906 21412
rect 434714 21400 434720 21412
rect 138900 21372 434720 21400
rect 138900 21360 138906 21372
rect 434714 21360 434720 21372
rect 434772 21360 434778 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 139394 20652 139400 20664
rect 3568 20624 139400 20652
rect 3568 20612 3574 20624
rect 139394 20612 139400 20624
rect 139452 20612 139458 20664
rect 180702 20612 180708 20664
rect 180760 20652 180766 20664
rect 580166 20652 580172 20664
rect 180760 20624 580172 20652
rect 180760 20612 180766 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 160002 18640 160008 18692
rect 160060 18680 160066 18692
rect 361574 18680 361580 18692
rect 160060 18652 361580 18680
rect 160060 18640 160066 18652
rect 361574 18640 361580 18652
rect 361632 18640 361638 18692
rect 134610 18572 134616 18624
rect 134668 18612 134674 18624
rect 454034 18612 454040 18624
rect 134668 18584 454040 18612
rect 134668 18572 134674 18584
rect 454034 18572 454040 18584
rect 454092 18572 454098 18624
rect 153838 17212 153844 17264
rect 153896 17252 153902 17264
rect 465074 17252 465080 17264
rect 153896 17224 465080 17252
rect 153896 17212 153902 17224
rect 465074 17212 465080 17224
rect 465132 17212 465138 17264
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 131206 16572 131212 16584
rect 3568 16544 131212 16572
rect 3568 16532 3574 16544
rect 131206 16532 131212 16544
rect 131264 16532 131270 16584
rect 165430 16532 165436 16584
rect 165488 16572 165494 16584
rect 580166 16572 580172 16584
rect 165488 16544 580172 16572
rect 165488 16532 165494 16544
rect 580166 16532 580172 16544
rect 580224 16532 580230 16584
rect 151078 14492 151084 14544
rect 151136 14532 151142 14544
rect 316402 14532 316408 14544
rect 151136 14504 316408 14532
rect 151136 14492 151142 14504
rect 316402 14492 316408 14504
rect 316460 14492 316466 14544
rect 166902 14424 166908 14476
rect 166960 14464 166966 14476
rect 549530 14464 549536 14476
rect 166960 14436 549536 14464
rect 166960 14424 166966 14436
rect 549530 14424 549536 14436
rect 549588 14424 549594 14476
rect 142890 13064 142896 13116
rect 142948 13104 142954 13116
rect 477218 13104 477224 13116
rect 142948 13076 477224 13104
rect 142948 13064 142954 13076
rect 477218 13064 477224 13076
rect 477276 13064 477282 13116
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 130378 12424 130384 12436
rect 3108 12396 130384 12424
rect 3108 12384 3114 12396
rect 130378 12384 130384 12396
rect 130436 12384 130442 12436
rect 182082 12384 182088 12436
rect 182140 12424 182146 12436
rect 580166 12424 580172 12436
rect 182140 12396 580172 12424
rect 182140 12384 182146 12396
rect 580166 12384 580172 12396
rect 580224 12384 580230 12436
rect 137186 10344 137192 10396
rect 137244 10384 137250 10396
rect 176010 10384 176016 10396
rect 137244 10356 176016 10384
rect 137244 10344 137250 10356
rect 176010 10344 176016 10356
rect 176068 10344 176074 10396
rect 142798 10276 142804 10328
rect 142856 10316 142862 10328
rect 418798 10316 418804 10328
rect 142856 10288 418804 10316
rect 142856 10276 142862 10288
rect 418798 10276 418804 10288
rect 418856 10276 418862 10328
rect 160370 9052 160376 9104
rect 160428 9092 160434 9104
rect 175918 9092 175924 9104
rect 160428 9064 175924 9092
rect 160428 9052 160434 9064
rect 175918 9052 175924 9064
rect 175976 9052 175982 9104
rect 145558 8984 145564 9036
rect 145616 9024 145622 9036
rect 340046 9024 340052 9036
rect 145616 8996 340052 9024
rect 145616 8984 145622 8996
rect 340046 8984 340052 8996
rect 340104 8984 340110 9036
rect 134518 8916 134524 8968
rect 134576 8956 134582 8968
rect 530670 8956 530676 8968
rect 134576 8928 530676 8956
rect 134576 8916 134582 8928
rect 530670 8916 530676 8928
rect 530728 8916 530734 8968
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 13078 8276 13084 8288
rect 3016 8248 13084 8276
rect 3016 8236 3022 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 152458 8236 152464 8288
rect 152516 8276 152522 8288
rect 580166 8276 580172 8288
rect 152516 8248 580172 8276
rect 152516 8236 152522 8248
rect 580166 8236 580172 8248
rect 580224 8236 580230 8288
rect 165522 7556 165528 7608
rect 165580 7596 165586 7608
rect 461762 7596 461768 7608
rect 165580 7568 461768 7596
rect 165580 7556 165586 7568
rect 461762 7556 461768 7568
rect 461820 7556 461826 7608
rect 162762 6128 162768 6180
rect 162820 6168 162826 6180
rect 473354 6168 473360 6180
rect 162820 6140 473360 6168
rect 162820 6128 162826 6140
rect 473354 6128 473360 6140
rect 473412 6128 473418 6180
rect 542998 5448 543004 5500
rect 543056 5488 543062 5500
rect 580166 5488 580172 5500
rect 543056 5460 580172 5488
rect 543056 5448 543062 5460
rect 580166 5448 580172 5460
rect 580224 5448 580230 5500
rect 152642 4836 152648 4888
rect 152700 4876 152706 4888
rect 171778 4876 171784 4888
rect 152700 4848 171784 4876
rect 152700 4836 152706 4848
rect 171778 4836 171784 4848
rect 171836 4836 171842 4888
rect 38010 4768 38016 4820
rect 38068 4808 38074 4820
rect 116578 4808 116584 4820
rect 38068 4780 116584 4808
rect 38068 4768 38074 4780
rect 116578 4768 116584 4780
rect 116636 4768 116642 4820
rect 158622 4768 158628 4820
rect 158680 4808 158686 4820
rect 542262 4808 542268 4820
rect 158680 4780 542268 4808
rect 158680 4768 158686 4780
rect 542262 4768 542268 4780
rect 542320 4768 542326 4820
rect 148778 4632 148784 4684
rect 148836 4672 148842 4684
rect 151906 4672 151912 4684
rect 148836 4644 151912 4672
rect 148836 4632 148842 4644
rect 151906 4632 151912 4644
rect 151964 4632 151970 4684
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 54478 4128 54484 4140
rect 3200 4100 54484 4128
rect 3200 4088 3206 4100
rect 54478 4088 54484 4100
rect 54536 4088 54542 4140
rect 34146 3680 34152 3732
rect 34204 3720 34210 3732
rect 36538 3720 36544 3732
rect 34204 3692 36544 3720
rect 34204 3680 34210 3692
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 174538 3612 174544 3664
rect 174596 3652 174602 3664
rect 186774 3652 186780 3664
rect 174596 3624 186780 3652
rect 174596 3612 174602 3624
rect 186774 3612 186780 3624
rect 186832 3612 186838 3664
rect 14 3544 20 3596
rect 72 3584 78 3596
rect 3326 3584 3332 3596
rect 72 3556 3332 3584
rect 72 3544 78 3556
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 91462 3544 91468 3596
rect 91520 3584 91526 3596
rect 93118 3584 93124 3596
rect 91520 3556 93124 3584
rect 91520 3544 91526 3556
rect 93118 3544 93124 3556
rect 93176 3544 93182 3596
rect 97810 3544 97816 3596
rect 97868 3584 97874 3596
rect 179046 3584 179052 3596
rect 97868 3556 179052 3584
rect 97868 3544 97874 3556
rect 179046 3544 179052 3556
rect 179104 3544 179110 3596
rect 242894 3544 242900 3596
rect 242952 3584 242958 3596
rect 244090 3584 244096 3596
rect 242952 3556 244096 3584
rect 242952 3544 242958 3556
rect 244090 3544 244096 3556
rect 244148 3544 244154 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 263410 3584 263416 3596
rect 262272 3556 263416 3584
rect 262272 3544 262278 3556
rect 263410 3544 263416 3556
rect 263468 3544 263474 3596
rect 265618 3544 265624 3596
rect 265676 3584 265682 3596
rect 267274 3584 267280 3596
rect 265676 3556 267280 3584
rect 265676 3544 265682 3556
rect 267274 3544 267280 3556
rect 267332 3544 267338 3596
rect 281534 3544 281540 3596
rect 281592 3584 281598 3596
rect 282730 3584 282736 3596
rect 281592 3556 282736 3584
rect 281592 3544 281598 3556
rect 282730 3544 282736 3556
rect 282788 3544 282794 3596
rect 357434 3544 357440 3596
rect 357492 3584 357498 3596
rect 358722 3584 358728 3596
rect 357492 3556 358728 3584
rect 357492 3544 357498 3556
rect 358722 3544 358728 3556
rect 358780 3544 358786 3596
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 4798 3516 4804 3528
rect 3292 3488 4804 3516
rect 3292 3476 3298 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 31018 3516 31024 3528
rect 30340 3488 31024 3516
rect 30340 3476 30346 3488
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 43438 3516 43444 3528
rect 41932 3488 43444 3516
rect 41932 3476 41938 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 48314 3476 48320 3528
rect 48372 3516 48378 3528
rect 49602 3516 49608 3528
rect 48372 3488 49608 3516
rect 48372 3476 48378 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 53466 3476 53472 3528
rect 53524 3516 53530 3528
rect 64138 3516 64144 3528
rect 53524 3488 64144 3516
rect 53524 3476 53530 3488
rect 64138 3476 64144 3488
rect 64196 3476 64202 3528
rect 72142 3476 72148 3528
rect 72200 3516 72206 3528
rect 72200 3488 135852 3516
rect 72200 3476 72206 3488
rect 64414 3408 64420 3460
rect 64472 3448 64478 3460
rect 135438 3448 135444 3460
rect 64472 3420 135444 3448
rect 64472 3408 64478 3420
rect 135438 3408 135444 3420
rect 135496 3408 135502 3460
rect 135824 3380 135852 3488
rect 135898 3476 135904 3528
rect 135956 3516 135962 3528
rect 141050 3516 141056 3528
rect 135956 3488 141056 3516
rect 135956 3476 135962 3488
rect 141050 3476 141056 3488
rect 141108 3476 141114 3528
rect 146938 3476 146944 3528
rect 146996 3516 147002 3528
rect 381906 3516 381912 3528
rect 146996 3488 381912 3516
rect 146996 3476 147002 3488
rect 381906 3476 381912 3488
rect 381964 3476 381970 3528
rect 395338 3476 395344 3528
rect 395396 3516 395402 3528
rect 416038 3516 416044 3528
rect 395396 3488 416044 3516
rect 395396 3476 395402 3488
rect 416038 3476 416044 3488
rect 416096 3476 416102 3528
rect 418798 3476 418804 3528
rect 418856 3516 418862 3528
rect 419902 3516 419908 3528
rect 418856 3488 419908 3516
rect 418856 3476 418862 3488
rect 419902 3476 419908 3488
rect 419960 3476 419966 3528
rect 442258 3476 442264 3528
rect 442316 3516 442322 3528
rect 443086 3516 443092 3528
rect 442316 3488 443092 3516
rect 442316 3476 442322 3488
rect 443086 3476 443092 3488
rect 443144 3476 443150 3528
rect 571334 3476 571340 3528
rect 571392 3516 571398 3528
rect 572530 3516 572536 3528
rect 571392 3488 572536 3516
rect 571392 3476 571398 3488
rect 572530 3476 572536 3488
rect 572588 3476 572594 3528
rect 138658 3408 138664 3460
rect 138716 3448 138722 3460
rect 557718 3448 557724 3460
rect 138716 3420 557724 3448
rect 138716 3408 138722 3420
rect 557718 3408 557724 3420
rect 557776 3408 557782 3460
rect 558178 3408 558184 3460
rect 558236 3448 558242 3460
rect 568666 3448 568672 3460
rect 558236 3420 568672 3448
rect 558236 3408 558242 3420
rect 568666 3408 568672 3420
rect 568724 3408 568730 3460
rect 139486 3380 139492 3392
rect 135824 3352 139492 3380
rect 139486 3340 139492 3352
rect 139544 3340 139550 3392
rect 211798 3000 211804 3052
rect 211856 3040 211862 3052
rect 213822 3040 213828 3052
rect 211856 3012 213828 3040
rect 211856 3000 211862 3012
rect 213822 3000 213828 3012
rect 213880 3000 213886 3052
rect 392578 3000 392584 3052
rect 392636 3040 392642 3052
rect 393498 3040 393504 3052
rect 392636 3012 393504 3040
rect 392636 3000 392642 3012
rect 393498 3000 393504 3012
rect 393556 3000 393562 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565446 3040 565452 3052
rect 563756 3012 565452 3040
rect 563756 3000 563762 3012
rect 565446 3000 565452 3012
rect 565504 3000 565510 3052
rect 376754 2592 376760 2644
rect 376812 2632 376818 2644
rect 378042 2632 378048 2644
rect 376812 2604 378048 2632
rect 376812 2592 376818 2604
rect 378042 2592 378048 2604
rect 378100 2592 378106 2644
rect 396074 2592 396080 2644
rect 396132 2632 396138 2644
rect 397362 2632 397368 2644
rect 396132 2604 397368 2632
rect 396132 2592 396138 2604
rect 397362 2592 397368 2604
rect 397420 2592 397426 2644
<< via1 >>
rect 49700 702992 49752 703044
rect 50896 702992 50948 703044
rect 69020 702992 69072 703044
rect 70216 702992 70268 703044
rect 309140 702992 309192 703044
rect 310428 702992 310480 703044
rect 328460 702992 328512 703044
rect 329748 702992 329800 703044
rect 347780 702992 347832 703044
rect 349068 702992 349120 703044
rect 358820 702992 358872 703044
rect 360016 702992 360068 703044
rect 378140 702992 378192 703044
rect 379336 702992 379388 703044
rect 576124 702448 576176 702500
rect 580172 702448 580224 702500
rect 3056 701020 3108 701072
rect 98644 701020 98696 701072
rect 184848 700612 184900 700664
rect 195980 700612 196032 700664
rect 188068 700544 188120 700596
rect 200120 700544 200172 700596
rect 66352 700476 66404 700528
rect 78036 700476 78088 700528
rect 115848 700476 115900 700528
rect 123668 700476 123720 700528
rect 177120 700476 177172 700528
rect 194692 700476 194744 700528
rect 19984 700408 20036 700460
rect 31024 700408 31076 700460
rect 77300 700408 77352 700460
rect 116032 700408 116084 700460
rect 169392 700408 169444 700460
rect 191840 700408 191892 700460
rect 194508 700408 194560 700460
rect 287888 700408 287940 700460
rect 16120 700340 16172 700392
rect 77944 700340 77996 700392
rect 117228 700340 117280 700392
rect 127532 700340 127584 700392
rect 165528 700340 165580 700392
rect 193220 700340 193272 700392
rect 199384 700340 199436 700392
rect 394792 700340 394844 700392
rect 548616 700340 548668 700392
rect 570604 700340 570656 700392
rect 31576 700272 31628 700324
rect 113180 700272 113232 700324
rect 121276 700272 121328 700324
rect 157800 700272 157852 700324
rect 189724 700272 189776 700324
rect 551284 700272 551336 700324
rect 556804 700272 556856 700324
rect 574468 700272 574520 700324
rect 180984 700068 181036 700120
rect 189448 700068 189500 700120
rect 115940 699796 115992 699848
rect 117964 699796 118016 699848
rect 119804 699660 119856 699712
rect 120724 699660 120776 699712
rect 199660 699660 199712 699712
rect 201500 699660 201552 699712
rect 220084 699660 220136 699712
rect 222844 699660 222896 699712
rect 224224 699660 224276 699712
rect 226708 699660 226760 699712
rect 242164 699660 242216 699712
rect 245384 699660 245436 699712
rect 269764 699660 269816 699712
rect 272432 699660 272484 699712
rect 278044 699660 278096 699712
rect 280160 699660 280212 699712
rect 323584 699660 323636 699712
rect 325884 699660 325936 699712
rect 374644 699660 374696 699712
rect 375472 699660 375524 699712
rect 395344 699660 395396 699712
rect 398656 699660 398708 699712
rect 400864 699660 400916 699712
rect 402520 699660 402572 699712
rect 445024 699660 445076 699712
rect 448244 699660 448296 699712
rect 449164 699660 449216 699712
rect 452108 699660 452160 699712
rect 472624 699660 472676 699712
rect 474648 699660 474700 699712
rect 494704 699660 494756 699712
rect 497832 699660 497884 699712
rect 498844 699660 498896 699712
rect 501696 699660 501748 699712
rect 502984 699660 503036 699712
rect 505560 699660 505612 699712
rect 552664 699660 552716 699712
rect 555148 699660 555200 699712
rect 570604 698300 570656 698352
rect 580172 698300 580224 698352
rect 144920 697552 144972 697604
rect 146208 697552 146260 697604
rect 492680 697552 492732 697604
rect 493968 697552 494020 697604
rect 512000 697552 512052 697604
rect 513288 697552 513340 697604
rect 544384 694152 544436 694204
rect 580172 694152 580224 694204
rect 3148 692792 3200 692844
rect 88984 692792 89036 692844
rect 3424 688644 3476 688696
rect 89076 688644 89128 688696
rect 548524 685856 548576 685908
rect 579804 685856 579856 685908
rect 3148 684496 3200 684548
rect 181444 684496 181496 684548
rect 3424 680348 3476 680400
rect 94504 680348 94556 680400
rect 576216 677560 576268 677612
rect 580172 677560 580224 677612
rect 3240 672052 3292 672104
rect 105544 672052 105596 672104
rect 556896 669332 556948 669384
rect 580172 669332 580224 669384
rect 3424 667904 3476 667956
rect 84844 667904 84896 667956
rect 202144 665184 202196 665236
rect 580172 665184 580224 665236
rect 3240 663756 3292 663808
rect 111892 663756 111944 663808
rect 3424 661036 3476 661088
rect 80704 661036 80756 661088
rect 3056 652740 3108 652792
rect 111064 652740 111116 652792
rect 196624 648592 196676 648644
rect 579988 648592 580040 648644
rect 3424 644444 3476 644496
rect 98736 644444 98788 644496
rect 566464 644444 566516 644496
rect 580172 644444 580224 644496
rect 567844 633428 567896 633480
rect 580172 633428 580224 633480
rect 552756 629280 552808 629332
rect 580172 629280 580224 629332
rect 3424 627920 3476 627972
rect 95884 627920 95936 627972
rect 577504 625404 577556 625456
rect 580540 625404 580592 625456
rect 3240 623772 3292 623824
rect 128360 623772 128412 623824
rect 3424 619624 3476 619676
rect 106924 619624 106976 619676
rect 3240 615476 3292 615528
rect 98828 615476 98880 615528
rect 3424 612756 3476 612808
rect 97264 612756 97316 612808
rect 3424 608608 3476 608660
rect 125692 608608 125744 608660
rect 565084 608608 565136 608660
rect 580172 608608 580224 608660
rect 3424 604460 3476 604512
rect 102784 604460 102836 604512
rect 3424 600312 3476 600364
rect 86224 600312 86276 600364
rect 3424 596164 3476 596216
rect 101404 596164 101456 596216
rect 567936 596164 567988 596216
rect 580172 596164 580224 596216
rect 198004 592016 198056 592068
rect 580172 592016 580224 592068
rect 3424 587868 3476 587920
rect 95976 587868 96028 587920
rect 3424 583720 3476 583772
rect 90364 583720 90416 583772
rect 574744 583720 574796 583772
rect 580172 583720 580224 583772
rect 3424 579640 3476 579692
rect 100024 579640 100076 579692
rect 3240 575492 3292 575544
rect 102876 575492 102928 575544
rect 566648 572704 566700 572756
rect 580172 572704 580224 572756
rect 3424 571344 3476 571396
rect 90456 571344 90508 571396
rect 544476 568556 544528 568608
rect 579712 568556 579764 568608
rect 3240 567196 3292 567248
rect 91744 567196 91796 567248
rect 3424 564408 3476 564460
rect 7564 564408 7616 564460
rect 571984 564408 572036 564460
rect 580172 564408 580224 564460
rect 3424 560260 3476 560312
rect 93124 560260 93176 560312
rect 200764 560260 200816 560312
rect 579620 560260 579672 560312
rect 3424 556180 3476 556232
rect 110420 556180 110472 556232
rect 3424 552032 3476 552084
rect 112444 552032 112496 552084
rect 3240 547884 3292 547936
rect 107016 547884 107068 547936
rect 193864 547884 193916 547936
rect 580080 547884 580132 547936
rect 3332 543736 3384 543788
rect 61384 543736 61436 543788
rect 554044 543736 554096 543788
rect 580172 543736 580224 543788
rect 3424 539588 3476 539640
rect 104164 539588 104216 539640
rect 570696 539588 570748 539640
rect 579712 539588 579764 539640
rect 192484 535440 192536 535492
rect 580172 535440 580224 535492
rect 3240 531292 3292 531344
rect 94596 531292 94648 531344
rect 3424 527144 3476 527196
rect 10324 527144 10376 527196
rect 560944 527144 560996 527196
rect 580172 527144 580224 527196
rect 3240 522996 3292 523048
rect 86316 522996 86368 523048
rect 562324 522996 562376 523048
rect 580172 522996 580224 523048
rect 3424 520276 3476 520328
rect 121460 520276 121512 520328
rect 574836 520276 574888 520328
rect 579712 520276 579764 520328
rect 3424 516128 3476 516180
rect 102968 516128 103020 516180
rect 573364 516128 573416 516180
rect 580172 516128 580224 516180
rect 3424 511980 3476 512032
rect 96344 511980 96396 512032
rect 566556 511980 566608 512032
rect 579620 511980 579672 512032
rect 3424 507832 3476 507884
rect 109684 507832 109736 507884
rect 558184 507832 558236 507884
rect 580172 507832 580224 507884
rect 3240 503684 3292 503736
rect 120816 503684 120868 503736
rect 192576 503684 192628 503736
rect 580080 503684 580132 503736
rect 3332 499536 3384 499588
rect 97356 499536 97408 499588
rect 576308 499536 576360 499588
rect 580172 499536 580224 499588
rect 2872 495456 2924 495508
rect 93216 495456 93268 495508
rect 558276 495456 558328 495508
rect 580172 495456 580224 495508
rect 3424 491308 3476 491360
rect 109776 491308 109828 491360
rect 3424 487160 3476 487212
rect 14464 487160 14516 487212
rect 569224 487160 569276 487212
rect 580172 487160 580224 487212
rect 3516 483012 3568 483064
rect 17224 483012 17276 483064
rect 182180 483012 182232 483064
rect 580172 483012 580224 483064
rect 3424 478864 3476 478916
rect 91836 478864 91888 478916
rect 563704 478864 563756 478916
rect 580172 478864 580224 478916
rect 3240 474716 3292 474768
rect 120080 474716 120132 474768
rect 561036 474716 561088 474768
rect 580172 474716 580224 474768
rect 3424 471996 3476 472048
rect 107200 471996 107252 472048
rect 561128 471996 561180 472048
rect 580172 471996 580224 472048
rect 3424 467848 3476 467900
rect 131120 467848 131172 467900
rect 563796 467848 563848 467900
rect 580172 467848 580224 467900
rect 3424 463700 3476 463752
rect 107108 463700 107160 463752
rect 562416 463700 562468 463752
rect 580172 463700 580224 463752
rect 3424 459552 3476 459604
rect 100116 459552 100168 459604
rect 552848 459552 552900 459604
rect 580172 459552 580224 459604
rect 3240 455404 3292 455456
rect 94688 455404 94740 455456
rect 558368 455404 558420 455456
rect 580080 455404 580132 455456
rect 3332 451256 3384 451308
rect 103612 451256 103664 451308
rect 124864 451256 124916 451308
rect 580172 451256 580224 451308
rect 572076 447108 572128 447160
rect 579712 447108 579764 447160
rect 3424 442960 3476 443012
rect 86408 442960 86460 443012
rect 561220 442960 561272 443012
rect 580172 442960 580224 443012
rect 570788 434732 570840 434784
rect 580172 434732 580224 434784
rect 3516 430584 3568 430636
rect 89168 430584 89220 430636
rect 568028 430584 568080 430636
rect 580172 430584 580224 430636
rect 2872 426436 2924 426488
rect 103060 426436 103112 426488
rect 563888 426436 563940 426488
rect 580172 426436 580224 426488
rect 574928 423648 574980 423700
rect 580172 423648 580224 423700
rect 2964 422288 3016 422340
rect 98920 422288 98972 422340
rect 3516 419500 3568 419552
rect 103152 419500 103204 419552
rect 191748 419500 191800 419552
rect 580172 419500 580224 419552
rect 3516 415420 3568 415472
rect 108304 415420 108356 415472
rect 210424 415420 210476 415472
rect 580172 415420 580224 415472
rect 3516 411272 3568 411324
rect 90548 411272 90600 411324
rect 575112 411272 575164 411324
rect 579988 411272 580040 411324
rect 3516 407124 3568 407176
rect 93308 407124 93360 407176
rect 124220 407124 124272 407176
rect 580172 407124 580224 407176
rect 3332 402976 3384 403028
rect 96160 402976 96212 403028
rect 565176 402976 565228 403028
rect 580172 402976 580224 403028
rect 179420 398828 179472 398880
rect 579712 398828 579764 398880
rect 576400 394680 576452 394732
rect 580172 394680 580224 394732
rect 3516 390532 3568 390584
rect 118700 390532 118752 390584
rect 572168 390532 572220 390584
rect 580172 390532 580224 390584
rect 3516 386384 3568 386436
rect 100208 386384 100260 386436
rect 189816 386384 189868 386436
rect 580172 386384 580224 386436
rect 2872 378156 2924 378208
rect 89260 378156 89312 378208
rect 184940 375368 184992 375420
rect 580172 375368 580224 375420
rect 2964 374008 3016 374060
rect 108396 374008 108448 374060
rect 555424 371220 555476 371272
rect 579804 371220 579856 371272
rect 3056 369860 3108 369912
rect 111156 369860 111208 369912
rect 189908 367072 189960 367124
rect 580172 367072 580224 367124
rect 3056 361564 3108 361616
rect 97448 361564 97500 361616
rect 3332 358776 3384 358828
rect 105636 358776 105688 358828
rect 566740 358776 566792 358828
rect 580172 358776 580224 358828
rect 3332 354696 3384 354748
rect 100300 354696 100352 354748
rect 178040 354696 178092 354748
rect 580172 354696 580224 354748
rect 3516 350548 3568 350600
rect 104256 350548 104308 350600
rect 206284 350548 206336 350600
rect 580172 350548 580224 350600
rect 3332 346400 3384 346452
rect 75184 346400 75236 346452
rect 569316 346400 569368 346452
rect 580172 346400 580224 346452
rect 3516 342252 3568 342304
rect 104900 342252 104952 342304
rect 563980 342252 564032 342304
rect 579712 342252 579764 342304
rect 3516 338104 3568 338156
rect 108488 338104 108540 338156
rect 577596 338104 577648 338156
rect 579620 338104 579672 338156
rect 572260 331236 572312 331288
rect 579712 331236 579764 331288
rect 2964 329808 3016 329860
rect 109868 329808 109920 329860
rect 3056 321580 3108 321632
rect 94780 321580 94832 321632
rect 577688 318792 577740 318844
rect 579712 318792 579764 318844
rect 3516 317432 3568 317484
rect 94872 317432 94924 317484
rect 575020 314644 575072 314696
rect 579620 314644 579672 314696
rect 3056 313284 3108 313336
rect 126980 313284 127032 313336
rect 558460 310496 558512 310548
rect 580172 310496 580224 310548
rect 3148 309136 3200 309188
rect 108580 309136 108632 309188
rect 564072 306348 564124 306400
rect 580172 306348 580224 306400
rect 3240 304988 3292 305040
rect 105728 304988 105780 305040
rect 569408 302200 569460 302252
rect 580172 302200 580224 302252
rect 3148 300840 3200 300892
rect 118792 300840 118844 300892
rect 3332 298120 3384 298172
rect 118056 298120 118108 298172
rect 3516 293972 3568 294024
rect 101496 293972 101548 294024
rect 170404 293972 170456 294024
rect 580172 293972 580224 294024
rect 3516 289824 3568 289876
rect 120264 289824 120316 289876
rect 558552 289824 558604 289876
rect 579988 289824 580040 289876
rect 2872 285676 2924 285728
rect 108672 285676 108724 285728
rect 572352 285676 572404 285728
rect 579988 285676 580040 285728
rect 555516 282888 555568 282940
rect 580172 282888 580224 282940
rect 2964 281528 3016 281580
rect 102692 281528 102744 281580
rect 561312 278740 561364 278792
rect 580172 278740 580224 278792
rect 122932 277992 122984 278044
rect 498844 277992 498896 278044
rect 3056 277380 3108 277432
rect 97816 277380 97868 277432
rect 195244 276632 195296 276684
rect 524420 276632 524472 276684
rect 169760 276020 169812 276072
rect 195244 276020 195296 276072
rect 566832 274660 566884 274712
rect 580172 274660 580224 274712
rect 147680 273912 147732 273964
rect 218060 273912 218112 273964
rect 3516 273232 3568 273284
rect 99932 273232 99984 273284
rect 191656 272484 191708 272536
rect 206284 272484 206336 272536
rect 155960 271872 156012 271924
rect 190460 271872 190512 271924
rect 191656 271872 191708 271924
rect 149152 271192 149204 271244
rect 202144 271192 202196 271244
rect 17224 271124 17276 271176
rect 110512 271124 110564 271176
rect 142804 271124 142856 271176
rect 230480 271124 230532 271176
rect 110512 270512 110564 270564
rect 111708 270512 111760 270564
rect 133972 270512 134024 270564
rect 577872 270512 577924 270564
rect 579712 270512 579764 270564
rect 132592 269764 132644 269816
rect 200764 269764 200816 269816
rect 3056 269084 3108 269136
rect 183652 269084 183704 269136
rect 10324 268404 10376 268456
rect 160100 268404 160152 268456
rect 145012 268336 145064 268388
rect 472624 268336 472676 268388
rect 111064 267724 111116 267776
rect 114468 267724 114520 267776
rect 139492 267724 139544 267776
rect 144828 267044 144880 267096
rect 170404 267044 170456 267096
rect 7564 266976 7616 267028
rect 167460 266976 167512 267028
rect 196992 266636 197044 266688
rect 198004 266636 198056 266688
rect 169760 266432 169812 266484
rect 198740 266432 198792 266484
rect 163964 266364 164016 266416
rect 196992 266364 197044 266416
rect 579620 266364 579672 266416
rect 189080 265956 189132 266008
rect 210424 265956 210476 266008
rect 161480 265888 161532 265940
rect 190000 265888 190052 265940
rect 153200 265820 153252 265872
rect 197360 265820 197412 265872
rect 133880 265752 133932 265804
rect 189632 265752 189684 265804
rect 136548 265684 136600 265736
rect 193864 265684 193916 265736
rect 148048 265616 148100 265668
rect 492680 265616 492732 265668
rect 3148 264936 3200 264988
rect 106832 264936 106884 264988
rect 118148 264936 118200 264988
rect 151912 264936 151964 264988
rect 154488 264936 154540 264988
rect 189080 264936 189132 264988
rect 189540 264936 189592 264988
rect 146208 264392 146260 264444
rect 192576 264392 192628 264444
rect 75184 264324 75236 264376
rect 158720 264324 158772 264376
rect 14464 264256 14516 264308
rect 158352 264256 158404 264308
rect 149244 264188 149296 264240
rect 150348 264188 150400 264240
rect 400864 264188 400916 264240
rect 115756 263984 115808 264036
rect 124864 263984 124916 264036
rect 125232 263984 125284 264036
rect 117136 263916 117188 263968
rect 126980 263916 127032 263968
rect 127716 263916 127768 263968
rect 114192 263848 114244 263900
rect 132592 263848 132644 263900
rect 133512 263848 133564 263900
rect 118516 263780 118568 263832
rect 145380 263780 145432 263832
rect 146208 263780 146260 263832
rect 115664 263712 115716 263764
rect 142620 263712 142672 263764
rect 166724 263712 166776 263764
rect 119988 263644 120040 263696
rect 149244 263644 149296 263696
rect 198924 263644 198976 263696
rect 112904 263576 112956 263628
rect 143724 263576 143776 263628
rect 144828 263576 144880 263628
rect 158720 263576 158772 263628
rect 159456 263576 159508 263628
rect 193588 263576 193640 263628
rect 132132 263508 132184 263560
rect 470600 263508 470652 263560
rect 23480 263440 23532 263492
rect 166724 263440 166776 263492
rect 57980 263372 58032 263424
rect 161940 263372 161992 263424
rect 69020 263304 69072 263356
rect 171600 263304 171652 263356
rect 157248 263100 157300 263152
rect 190828 263100 190880 263152
rect 267740 263100 267792 263152
rect 130016 263032 130068 263084
rect 276020 263032 276072 263084
rect 196256 262964 196308 263016
rect 347780 262964 347832 263016
rect 111064 262896 111116 262948
rect 126980 262896 127032 262948
rect 140780 262896 140832 262948
rect 299480 262896 299532 262948
rect 121552 262828 121604 262880
rect 138480 262828 138532 262880
rect 164792 262828 164844 262880
rect 194600 262828 194652 262880
rect 197636 262828 197688 262880
rect 119804 262760 119856 262812
rect 152556 262760 152608 262812
rect 155684 262760 155736 262812
rect 190644 262760 190696 262812
rect 119620 262692 119672 262744
rect 153384 262692 153436 262744
rect 170588 262692 170640 262744
rect 191104 262692 191156 262744
rect 119896 262624 119948 262676
rect 137652 262624 137704 262676
rect 174728 262624 174780 262676
rect 197544 262624 197596 262676
rect 116308 262556 116360 262608
rect 140136 262556 140188 262608
rect 173808 262556 173860 262608
rect 199108 262556 199160 262608
rect 477500 262828 477552 262880
rect 112996 262488 113048 262540
rect 136824 262488 136876 262540
rect 165528 262488 165580 262540
rect 192852 262488 192904 262540
rect 115572 262420 115624 262472
rect 141792 262420 141844 262472
rect 160652 262420 160704 262472
rect 193312 262420 193364 262472
rect 114284 262352 114336 262404
rect 140780 262352 140832 262404
rect 158168 262352 158220 262404
rect 190736 262352 190788 262404
rect 118240 262284 118292 262336
rect 130200 262284 130252 262336
rect 177948 262284 178000 262336
rect 179420 262284 179472 262336
rect 181352 262284 181404 262336
rect 196256 262284 196308 262336
rect 134892 262216 134944 262268
rect 135996 262216 136048 262268
rect 173072 262216 173124 262268
rect 193404 262216 193456 262268
rect 577780 262216 577832 262268
rect 580264 262216 580316 262268
rect 162768 260992 162820 261044
rect 3056 260924 3108 260976
rect 109960 260924 110012 260976
rect 111340 260924 111392 260976
rect 144828 260924 144880 260976
rect 192576 260924 192628 260976
rect 7564 260856 7616 260908
rect 176660 260856 176712 260908
rect 192392 260856 192444 260908
rect 193496 260856 193548 260908
rect 498844 260856 498896 260908
rect 118424 260788 118476 260840
rect 122840 260788 122892 260840
rect 129740 260788 129792 260840
rect 129924 260788 129976 260840
rect 132684 260788 132736 260840
rect 161204 260312 161256 260364
rect 194968 260312 195020 260364
rect 113824 260244 113876 260296
rect 124404 260244 124456 260296
rect 158352 260244 158404 260296
rect 193772 260244 193824 260296
rect 119712 260176 119764 260228
rect 144920 260176 144972 260228
rect 145012 260176 145064 260228
rect 146254 260176 146306 260228
rect 147680 260176 147732 260228
rect 148738 260176 148790 260228
rect 149060 260176 149112 260228
rect 190552 260176 190604 260228
rect 115480 260108 115532 260160
rect 129740 260108 129792 260160
rect 142160 260108 142212 260160
rect 192300 260108 192352 260160
rect 120172 260040 120224 260092
rect 121368 260040 121420 260092
rect 160100 260040 160152 260092
rect 161158 260040 161210 260092
rect 178040 260040 178092 260092
rect 179374 260040 179426 260092
rect 115204 259972 115256 260024
rect 126060 259972 126112 260024
rect 180340 259972 180392 260024
rect 192024 260040 192076 260092
rect 184664 259972 184716 260024
rect 196440 259972 196492 260024
rect 114008 259904 114060 259956
rect 123208 259904 123260 259956
rect 123576 259904 123628 259956
rect 178868 259904 178920 259956
rect 197728 259904 197780 259956
rect 116676 259836 116728 259888
rect 128452 259836 128504 259888
rect 179512 259836 179564 259888
rect 197912 259836 197964 259888
rect 112536 259768 112588 259820
rect 131120 259768 131172 259820
rect 167920 259768 167972 259820
rect 192208 259768 192260 259820
rect 115388 259700 115440 259752
rect 145012 259700 145064 259752
rect 172244 259700 172296 259752
rect 197820 259700 197872 259752
rect 116768 259632 116820 259684
rect 147680 259632 147732 259684
rect 166448 259632 166500 259684
rect 197084 259632 197136 259684
rect 113916 259564 113968 259616
rect 146760 259564 146812 259616
rect 162308 259564 162360 259616
rect 195244 259564 195296 259616
rect 116584 259496 116636 259548
rect 149152 259496 149204 259548
rect 175372 259496 175424 259548
rect 192116 259496 192168 259548
rect 117872 259428 117924 259480
rect 150900 259428 150952 259480
rect 176384 259428 176436 259480
rect 195060 259428 195112 259480
rect 3240 256708 3292 256760
rect 117320 256708 117372 256760
rect 191656 253920 191708 253972
rect 579804 253920 579856 253972
rect 120080 253172 120132 253224
rect 120356 253172 120408 253224
rect 3148 252560 3200 252612
rect 119344 252560 119396 252612
rect 192576 251132 192628 251184
rect 579988 251132 580040 251184
rect 191196 241476 191248 241528
rect 580172 241476 580224 241528
rect 3332 240116 3384 240168
rect 119436 240116 119488 240168
rect 498844 238688 498896 238740
rect 580172 238688 580224 238740
rect 3332 229100 3384 229152
rect 120908 229100 120960 229152
rect 190092 224952 190144 225004
rect 579988 224952 580040 225004
rect 3056 220804 3108 220856
rect 119528 220804 119580 220856
rect 3148 208360 3200 208412
rect 120540 208360 120592 208412
rect 190552 204892 190604 204944
rect 190920 204892 190972 204944
rect 96068 201492 96120 201544
rect 118700 201492 118752 201544
rect 118976 201492 119028 201544
rect 191472 201492 191524 201544
rect 191748 201492 191800 201544
rect 204260 201492 204312 201544
rect 115940 201424 115992 201476
rect 117044 201424 117096 201476
rect 3608 200812 3660 200864
rect 95148 200812 95200 200864
rect 96252 200812 96304 200864
rect 117320 200812 117372 200864
rect 3516 200744 3568 200796
rect 96436 200744 96488 200796
rect 109960 200744 110012 200796
rect 104532 200472 104584 200524
rect 113180 200472 113232 200524
rect 204352 200812 204404 200864
rect 252560 200812 252612 200864
rect 121184 200744 121236 200796
rect 125554 200676 125606 200728
rect 125692 200676 125744 200728
rect 119528 200608 119580 200660
rect 119344 200540 119396 200592
rect 132132 200540 132184 200592
rect 121184 200472 121236 200524
rect 124404 200472 124456 200524
rect 131764 200472 131816 200524
rect 131856 200472 131908 200524
rect 104440 200404 104492 200456
rect 118792 200404 118844 200456
rect 120540 200404 120592 200456
rect 121000 200404 121052 200456
rect 97540 200336 97592 200388
rect 115940 200336 115992 200388
rect 94964 200268 95016 200320
rect 120264 200268 120316 200320
rect 123208 200268 123260 200320
rect 96436 200200 96488 200252
rect 132132 200268 132184 200320
rect 132040 200200 132092 200252
rect 95148 200132 95200 200184
rect 131856 200132 131908 200184
rect 131948 200132 132000 200184
rect 129740 199996 129792 200048
rect 131856 199928 131908 199980
rect 121000 199792 121052 199844
rect 132224 199860 132276 199912
rect 132638 199860 132690 199912
rect 127900 199792 127952 199844
rect 119344 199724 119396 199776
rect 131856 199792 131908 199844
rect 133006 199860 133058 199912
rect 133098 199860 133150 199912
rect 132730 199792 132782 199844
rect 84200 199520 84252 199572
rect 128452 199520 128504 199572
rect 129648 199520 129700 199572
rect 133144 199724 133196 199776
rect 131764 199656 131816 199708
rect 133788 199656 133840 199708
rect 134018 199860 134070 199912
rect 134110 199860 134162 199912
rect 134570 199860 134622 199912
rect 134938 199860 134990 199912
rect 134156 199724 134208 199776
rect 134064 199656 134116 199708
rect 133696 199588 133748 199640
rect 134524 199588 134576 199640
rect 134892 199588 134944 199640
rect 131672 199520 131724 199572
rect 131856 199520 131908 199572
rect 133604 199520 133656 199572
rect 133788 199520 133840 199572
rect 134340 199520 134392 199572
rect 135398 199860 135450 199912
rect 135766 199860 135818 199912
rect 135720 199588 135772 199640
rect 135352 199520 135404 199572
rect 136042 199860 136094 199912
rect 136134 199860 136186 199912
rect 136226 199860 136278 199912
rect 136410 199860 136462 199912
rect 136088 199724 136140 199776
rect 136180 199724 136232 199776
rect 136456 199656 136508 199708
rect 136364 199588 136416 199640
rect 137238 199860 137290 199912
rect 136686 199792 136738 199844
rect 137146 199792 137198 199844
rect 137330 199792 137382 199844
rect 137192 199656 137244 199708
rect 137284 199656 137336 199708
rect 137606 199860 137658 199912
rect 137698 199860 137750 199912
rect 137790 199860 137842 199912
rect 137652 199724 137704 199776
rect 137744 199656 137796 199708
rect 137974 199860 138026 199912
rect 138710 199860 138762 199912
rect 138802 199860 138854 199912
rect 138894 199860 138946 199912
rect 139170 199860 139222 199912
rect 139446 199860 139498 199912
rect 137836 199588 137888 199640
rect 137468 199520 137520 199572
rect 138296 199520 138348 199572
rect 138480 199520 138532 199572
rect 138848 199724 138900 199776
rect 138848 199520 138900 199572
rect 139400 199724 139452 199776
rect 139722 199860 139774 199912
rect 139906 199860 139958 199912
rect 140458 199860 140510 199912
rect 140642 199860 140694 199912
rect 140826 199860 140878 199912
rect 141102 199860 141154 199912
rect 141194 199860 141246 199912
rect 141286 199860 141338 199912
rect 141378 199860 141430 199912
rect 139124 199588 139176 199640
rect 139492 199588 139544 199640
rect 139676 199588 139728 199640
rect 139860 199588 139912 199640
rect 140320 199588 140372 199640
rect 46940 199452 46992 199504
rect 138940 199452 138992 199504
rect 4068 199384 4120 199436
rect 121276 199316 121328 199368
rect 140044 199316 140096 199368
rect 141240 199724 141292 199776
rect 141148 199656 141200 199708
rect 141332 199656 141384 199708
rect 140964 199588 141016 199640
rect 141056 199588 141108 199640
rect 141516 199588 141568 199640
rect 141930 199860 141982 199912
rect 142206 199860 142258 199912
rect 142298 199860 142350 199912
rect 142390 199860 142442 199912
rect 142574 199860 142626 199912
rect 142666 199860 142718 199912
rect 142758 199860 142810 199912
rect 142850 199860 142902 199912
rect 142160 199724 142212 199776
rect 142436 199724 142488 199776
rect 142620 199724 142672 199776
rect 142896 199724 142948 199776
rect 142252 199656 142304 199708
rect 142528 199656 142580 199708
rect 142712 199656 142764 199708
rect 143494 199860 143546 199912
rect 143770 199860 143822 199912
rect 144046 199860 144098 199912
rect 143080 199588 143132 199640
rect 142436 199520 142488 199572
rect 143724 199520 143776 199572
rect 144000 199520 144052 199572
rect 144322 199860 144374 199912
rect 144460 199588 144512 199640
rect 141056 199452 141108 199504
rect 142712 199452 142764 199504
rect 143448 199452 143500 199504
rect 144092 199452 144144 199504
rect 140596 199384 140648 199436
rect 140780 199384 140832 199436
rect 144690 199860 144742 199912
rect 144782 199860 144834 199912
rect 145058 199860 145110 199912
rect 145426 199860 145478 199912
rect 145518 199860 145570 199912
rect 145610 199860 145662 199912
rect 145886 199860 145938 199912
rect 144736 199656 144788 199708
rect 145242 199792 145294 199844
rect 144644 199520 144696 199572
rect 145012 199520 145064 199572
rect 144736 199452 144788 199504
rect 145472 199656 145524 199708
rect 145564 199656 145616 199708
rect 145380 199588 145432 199640
rect 146254 199860 146306 199912
rect 146346 199860 146398 199912
rect 146530 199860 146582 199912
rect 146806 199860 146858 199912
rect 146898 199860 146950 199912
rect 147174 199860 147226 199912
rect 147266 199860 147318 199912
rect 146622 199792 146674 199844
rect 146484 199656 146536 199708
rect 146668 199656 146720 199708
rect 146990 199792 147042 199844
rect 146944 199656 146996 199708
rect 146392 199588 146444 199640
rect 146760 199588 146812 199640
rect 146300 199520 146352 199572
rect 146576 199520 146628 199572
rect 147634 199860 147686 199912
rect 147726 199860 147778 199912
rect 147220 199588 147272 199640
rect 147496 199588 147548 199640
rect 107568 199248 107620 199300
rect 133604 199248 133656 199300
rect 135076 199248 135128 199300
rect 135628 199248 135680 199300
rect 138020 199248 138072 199300
rect 145656 199248 145708 199300
rect 129648 199180 129700 199232
rect 141424 199180 141476 199232
rect 145840 199316 145892 199368
rect 146576 199248 146628 199300
rect 147680 199656 147732 199708
rect 147910 199860 147962 199912
rect 148002 199860 148054 199912
rect 148094 199860 148146 199912
rect 147956 199724 148008 199776
rect 148278 199860 148330 199912
rect 148554 199860 148606 199912
rect 148646 199860 148698 199912
rect 148922 199860 148974 199912
rect 149106 199860 149158 199912
rect 148462 199792 148514 199844
rect 148232 199656 148284 199708
rect 147864 199588 147916 199640
rect 148140 199588 148192 199640
rect 148048 199520 148100 199572
rect 148830 199724 148882 199776
rect 148968 199724 149020 199776
rect 148784 199520 148836 199572
rect 147864 199452 147916 199504
rect 148876 199316 148928 199368
rect 149382 199860 149434 199912
rect 149428 199724 149480 199776
rect 149842 199860 149894 199912
rect 150026 199860 150078 199912
rect 150118 199860 150170 199912
rect 150210 199860 150262 199912
rect 150394 199860 150446 199912
rect 150578 199860 150630 199912
rect 150072 199724 150124 199776
rect 150348 199724 150400 199776
rect 150854 199860 150906 199912
rect 150762 199792 150814 199844
rect 150624 199724 150676 199776
rect 150164 199656 150216 199708
rect 149980 199588 150032 199640
rect 150256 199520 150308 199572
rect 150716 199520 150768 199572
rect 149796 199452 149848 199504
rect 151314 199860 151366 199912
rect 151406 199860 151458 199912
rect 151590 199860 151642 199912
rect 151130 199724 151182 199776
rect 151360 199724 151412 199776
rect 151682 199792 151734 199844
rect 151636 199656 151688 199708
rect 151544 199520 151596 199572
rect 150992 199452 151044 199504
rect 151176 199452 151228 199504
rect 151268 199452 151320 199504
rect 151728 199452 151780 199504
rect 150256 199180 150308 199232
rect 150440 199180 150492 199232
rect 151636 199316 151688 199368
rect 150808 199248 150860 199300
rect 152418 199860 152470 199912
rect 153154 199860 153206 199912
rect 153246 199860 153298 199912
rect 152050 199792 152102 199844
rect 152234 199792 152286 199844
rect 152602 199792 152654 199844
rect 152096 199588 152148 199640
rect 152464 199588 152516 199640
rect 152372 199452 152424 199504
rect 152786 199792 152838 199844
rect 152924 199656 152976 199708
rect 152832 199588 152884 199640
rect 153476 199520 153528 199572
rect 153890 199860 153942 199912
rect 153982 199860 154034 199912
rect 154074 199860 154126 199912
rect 154258 199860 154310 199912
rect 154028 199724 154080 199776
rect 153200 199384 153252 199436
rect 153384 199384 153436 199436
rect 153752 199384 153804 199436
rect 153844 199384 153896 199436
rect 120264 199112 120316 199164
rect 125692 199044 125744 199096
rect 135996 199044 136048 199096
rect 138940 199044 138992 199096
rect 142988 199044 143040 199096
rect 145196 199044 145248 199096
rect 150256 199044 150308 199096
rect 151912 199112 151964 199164
rect 153108 199180 153160 199232
rect 154212 199588 154264 199640
rect 154442 199860 154494 199912
rect 154626 199860 154678 199912
rect 154718 199860 154770 199912
rect 154810 199860 154862 199912
rect 154902 199860 154954 199912
rect 154994 199860 155046 199912
rect 155362 199860 155414 199912
rect 154488 199656 154540 199708
rect 154580 199656 154632 199708
rect 154672 199656 154724 199708
rect 154764 199656 154816 199708
rect 154856 199656 154908 199708
rect 154396 199588 154448 199640
rect 155638 199860 155690 199912
rect 155730 199860 155782 199912
rect 156098 199860 156150 199912
rect 156190 199860 156242 199912
rect 156282 199860 156334 199912
rect 156374 199860 156426 199912
rect 155500 199588 155552 199640
rect 155684 199724 155736 199776
rect 156236 199656 156288 199708
rect 156328 199656 156380 199708
rect 156650 199860 156702 199912
rect 156742 199860 156794 199912
rect 156834 199860 156886 199912
rect 157110 199860 157162 199912
rect 157386 199860 157438 199912
rect 155960 199588 156012 199640
rect 156144 199588 156196 199640
rect 156512 199588 156564 199640
rect 156926 199792 156978 199844
rect 156788 199724 156840 199776
rect 157064 199656 157116 199708
rect 156696 199588 156748 199640
rect 156972 199588 157024 199640
rect 157340 199588 157392 199640
rect 157754 199860 157806 199912
rect 157938 199860 157990 199912
rect 158030 199860 158082 199912
rect 158122 199860 158174 199912
rect 158076 199588 158128 199640
rect 156880 199520 156932 199572
rect 157616 199520 157668 199572
rect 157708 199520 157760 199572
rect 157892 199520 157944 199572
rect 155224 199452 155276 199504
rect 158398 199860 158450 199912
rect 158490 199860 158542 199912
rect 158674 199860 158726 199912
rect 159502 199860 159554 199912
rect 159778 199860 159830 199912
rect 159870 199860 159922 199912
rect 158352 199656 158404 199708
rect 158444 199656 158496 199708
rect 158628 199588 158680 199640
rect 158536 199520 158588 199572
rect 159824 199656 159876 199708
rect 160100 199588 160152 199640
rect 156236 199384 156288 199436
rect 157156 199384 157208 199436
rect 158812 199452 158864 199504
rect 160514 199860 160566 199912
rect 160698 199860 160750 199912
rect 160790 199860 160842 199912
rect 160330 199792 160382 199844
rect 160422 199724 160474 199776
rect 160284 199656 160336 199708
rect 160376 199588 160428 199640
rect 160468 199520 160520 199572
rect 160560 199452 160612 199504
rect 160974 199860 161026 199912
rect 160836 199588 160888 199640
rect 161158 199860 161210 199912
rect 161342 199860 161394 199912
rect 161434 199860 161486 199912
rect 161526 199860 161578 199912
rect 161618 199860 161670 199912
rect 161710 199860 161762 199912
rect 161894 199860 161946 199912
rect 161986 199860 162038 199912
rect 162078 199860 162130 199912
rect 162262 199860 162314 199912
rect 161296 199724 161348 199776
rect 161204 199656 161256 199708
rect 161572 199724 161624 199776
rect 161020 199520 161072 199572
rect 161388 199588 161440 199640
rect 160744 199384 160796 199436
rect 154948 199316 155000 199368
rect 157340 199316 157392 199368
rect 161756 199588 161808 199640
rect 162032 199588 162084 199640
rect 162492 199520 162544 199572
rect 161940 199452 161992 199504
rect 162216 199384 162268 199436
rect 162906 199860 162958 199912
rect 163090 199860 163142 199912
rect 163182 199860 163234 199912
rect 163274 199860 163326 199912
rect 163734 199860 163786 199912
rect 162768 199588 162820 199640
rect 163044 199588 163096 199640
rect 163228 199520 163280 199572
rect 163044 199452 163096 199504
rect 163780 199452 163832 199504
rect 164194 199860 164246 199912
rect 164102 199792 164154 199844
rect 164056 199656 164108 199708
rect 164148 199656 164200 199708
rect 163964 199452 164016 199504
rect 164240 199452 164292 199504
rect 164470 199860 164522 199912
rect 164654 199860 164706 199912
rect 164746 199860 164798 199912
rect 164838 199860 164890 199912
rect 164930 199860 164982 199912
rect 165114 199860 165166 199912
rect 164700 199520 164752 199572
rect 164516 199452 164568 199504
rect 164608 199452 164660 199504
rect 164884 199656 164936 199708
rect 165068 199588 165120 199640
rect 164884 199452 164936 199504
rect 165850 199860 165902 199912
rect 165942 199860 165994 199912
rect 166126 199860 166178 199912
rect 166310 199792 166362 199844
rect 166080 199724 166132 199776
rect 165988 199656 166040 199708
rect 166264 199656 166316 199708
rect 166678 199860 166730 199912
rect 166770 199860 166822 199912
rect 167138 199860 167190 199912
rect 167230 199860 167282 199912
rect 166724 199724 166776 199776
rect 167046 199792 167098 199844
rect 165252 199384 165304 199436
rect 165436 199316 165488 199368
rect 165896 199384 165948 199436
rect 167092 199656 167144 199708
rect 166632 199316 166684 199368
rect 580724 200744 580776 200796
rect 562324 200676 562376 200728
rect 177948 200608 178000 200660
rect 191748 200608 191800 200660
rect 167414 199860 167466 199912
rect 167782 199860 167834 199912
rect 167874 199860 167926 199912
rect 167966 199860 168018 199912
rect 168058 199860 168110 199912
rect 168150 199860 168202 199912
rect 168334 199860 168386 199912
rect 168426 199860 168478 199912
rect 167276 199520 167328 199572
rect 167644 199520 167696 199572
rect 168012 199520 168064 199572
rect 168104 199520 168156 199572
rect 167920 199452 167972 199504
rect 167184 199384 167236 199436
rect 168380 199656 168432 199708
rect 169070 199860 169122 199912
rect 169346 199860 169398 199912
rect 169300 199724 169352 199776
rect 168564 199588 168616 199640
rect 169116 199588 169168 199640
rect 169622 199860 169674 199912
rect 169622 199656 169674 199708
rect 169392 199520 169444 199572
rect 169806 199860 169858 199912
rect 169990 199860 170042 199912
rect 170082 199860 170134 199912
rect 170174 199860 170226 199912
rect 170450 199860 170502 199912
rect 170542 199860 170594 199912
rect 171002 199860 171054 199912
rect 171278 199860 171330 199912
rect 171370 199860 171422 199912
rect 171462 199860 171514 199912
rect 171830 199860 171882 199912
rect 171922 199860 171974 199912
rect 169944 199724 169996 199776
rect 170128 199724 170180 199776
rect 170496 199724 170548 199776
rect 170588 199724 170640 199776
rect 170956 199724 171008 199776
rect 170036 199656 170088 199708
rect 171416 199724 171468 199776
rect 171600 199520 171652 199572
rect 171968 199724 172020 199776
rect 172382 199860 172434 199912
rect 172566 199860 172618 199912
rect 172842 199860 172894 199912
rect 172934 199860 172986 199912
rect 173026 199860 173078 199912
rect 173210 199860 173262 199912
rect 173486 199860 173538 199912
rect 173670 199860 173722 199912
rect 178684 200404 178736 200456
rect 178776 200200 178828 200252
rect 194508 200268 194560 200320
rect 211436 200268 211488 200320
rect 190552 200200 190604 200252
rect 191656 200200 191708 200252
rect 215392 200200 215444 200252
rect 204352 200132 204404 200184
rect 178408 200064 178460 200116
rect 173946 199860 173998 199912
rect 174038 199860 174090 199912
rect 174130 199860 174182 199912
rect 174406 199860 174458 199912
rect 174590 199860 174642 199912
rect 174774 199860 174826 199912
rect 172198 199724 172250 199776
rect 172428 199656 172480 199708
rect 172796 199724 172848 199776
rect 172888 199656 172940 199708
rect 173164 199724 173216 199776
rect 172152 199588 172204 199640
rect 172612 199588 172664 199640
rect 172980 199588 173032 199640
rect 173992 199724 174044 199776
rect 173854 199656 173906 199708
rect 174452 199724 174504 199776
rect 174728 199724 174780 199776
rect 174636 199656 174688 199708
rect 173532 199588 173584 199640
rect 180524 199996 180576 200048
rect 174958 199860 175010 199912
rect 175050 199860 175102 199912
rect 175142 199860 175194 199912
rect 175234 199860 175286 199912
rect 175418 199860 175470 199912
rect 175694 199860 175746 199912
rect 176154 199860 176206 199912
rect 175096 199724 175148 199776
rect 175096 199588 175148 199640
rect 168472 199452 168524 199504
rect 169668 199452 169720 199504
rect 171232 199452 171284 199504
rect 172244 199520 172296 199572
rect 174268 199520 174320 199572
rect 174912 199520 174964 199572
rect 175004 199520 175056 199572
rect 175326 199724 175378 199776
rect 175372 199588 175424 199640
rect 175878 199792 175930 199844
rect 175740 199656 175792 199708
rect 175832 199656 175884 199708
rect 176522 199860 176574 199912
rect 176338 199792 176390 199844
rect 176292 199588 176344 199640
rect 176384 199588 176436 199640
rect 181812 199928 181864 199980
rect 176706 199860 176758 199912
rect 177166 199860 177218 199912
rect 177350 199860 177402 199912
rect 180432 199860 180484 199912
rect 178040 199792 178092 199844
rect 177672 199724 177724 199776
rect 188988 199724 189040 199776
rect 192484 199724 192536 199776
rect 182272 199656 182324 199708
rect 178960 199588 179012 199640
rect 302240 199588 302292 199640
rect 171784 199452 171836 199504
rect 184756 199520 184808 199572
rect 189816 199520 189868 199572
rect 176660 199452 176712 199504
rect 176936 199452 176988 199504
rect 184940 199452 184992 199504
rect 186228 199452 186280 199504
rect 199384 199520 199436 199572
rect 216680 199520 216732 199572
rect 427820 199520 427872 199572
rect 201408 199452 201460 199504
rect 412640 199452 412692 199504
rect 168656 199384 168708 199436
rect 170772 199384 170824 199436
rect 431960 199384 432012 199436
rect 167368 199316 167420 199368
rect 170312 199316 170364 199368
rect 182180 199316 182232 199368
rect 156236 199248 156288 199300
rect 156972 199248 157024 199300
rect 157248 199248 157300 199300
rect 291200 199248 291252 199300
rect 159640 199180 159692 199232
rect 216680 199180 216732 199232
rect 152740 199112 152792 199164
rect 154028 199112 154080 199164
rect 155500 199112 155552 199164
rect 190552 199112 190604 199164
rect 152648 199044 152700 199096
rect 154948 199044 155000 199096
rect 160100 199044 160152 199096
rect 184940 199044 184992 199096
rect 130384 198976 130436 199028
rect 147956 198976 148008 199028
rect 190092 198976 190144 199028
rect 117964 198908 118016 198960
rect 164056 198908 164108 198960
rect 164240 198908 164292 198960
rect 164792 198908 164844 198960
rect 120724 198840 120776 198892
rect 124312 198840 124364 198892
rect 125508 198840 125560 198892
rect 128912 198840 128964 198892
rect 133144 198840 133196 198892
rect 135904 198840 135956 198892
rect 140964 198840 141016 198892
rect 142712 198840 142764 198892
rect 145196 198840 145248 198892
rect 145656 198840 145708 198892
rect 157248 198840 157300 198892
rect 160836 198840 160888 198892
rect 163596 198840 163648 198892
rect 120908 198772 120960 198824
rect 175556 198908 175608 198960
rect 175832 198908 175884 198960
rect 176200 198908 176252 198960
rect 176568 198908 176620 198960
rect 178040 198908 178092 198960
rect 165436 198840 165488 198892
rect 166172 198840 166224 198892
rect 169208 198840 169260 198892
rect 120816 198704 120868 198756
rect 124772 198704 124824 198756
rect 125508 198704 125560 198756
rect 144552 198704 144604 198756
rect 120724 198636 120776 198688
rect 121184 198568 121236 198620
rect 126520 198636 126572 198688
rect 134524 198636 134576 198688
rect 136272 198636 136324 198688
rect 144000 198636 144052 198688
rect 97724 198500 97776 198552
rect 121276 198500 121328 198552
rect 138388 198568 138440 198620
rect 103428 198432 103480 198484
rect 129740 198432 129792 198484
rect 102048 198364 102100 198416
rect 126520 198364 126572 198416
rect 143080 198500 143132 198552
rect 146024 198500 146076 198552
rect 173440 198772 173492 198824
rect 173624 198772 173676 198824
rect 174636 198840 174688 198892
rect 177764 198840 177816 198892
rect 185400 198840 185452 198892
rect 178960 198772 179012 198824
rect 179512 198772 179564 198824
rect 151636 198704 151688 198756
rect 155224 198704 155276 198756
rect 150256 198636 150308 198688
rect 154856 198636 154908 198688
rect 150716 198568 150768 198620
rect 165436 198704 165488 198756
rect 167644 198704 167696 198756
rect 168380 198704 168432 198756
rect 165620 198636 165672 198688
rect 184848 198704 184900 198756
rect 189908 198704 189960 198756
rect 172980 198636 173032 198688
rect 174084 198636 174136 198688
rect 182272 198636 182324 198688
rect 200396 198636 200448 198688
rect 201408 198636 201460 198688
rect 163596 198568 163648 198620
rect 169852 198568 169904 198620
rect 175648 198568 175700 198620
rect 195980 198568 196032 198620
rect 159732 198500 159784 198552
rect 169208 198500 169260 198552
rect 171508 198500 171560 198552
rect 173072 198500 173124 198552
rect 177028 198500 177080 198552
rect 194508 198500 194560 198552
rect 134616 198432 134668 198484
rect 140872 198432 140924 198484
rect 142436 198432 142488 198484
rect 161112 198432 161164 198484
rect 161940 198432 161992 198484
rect 162860 198432 162912 198484
rect 166264 198432 166316 198484
rect 183560 198432 183612 198484
rect 136824 198364 136876 198416
rect 141516 198364 141568 198416
rect 147956 198364 148008 198416
rect 155868 198364 155920 198416
rect 165436 198364 165488 198416
rect 165896 198364 165948 198416
rect 169208 198364 169260 198416
rect 170588 198364 170640 198416
rect 177672 198364 177724 198416
rect 100668 198296 100720 198348
rect 133696 198296 133748 198348
rect 144092 198296 144144 198348
rect 145104 198296 145156 198348
rect 156880 198296 156932 198348
rect 165712 198296 165764 198348
rect 168472 198296 168524 198348
rect 189264 198296 189316 198348
rect 101956 198228 102008 198280
rect 134432 198228 134484 198280
rect 100392 198160 100444 198212
rect 126152 198160 126204 198212
rect 148048 198228 148100 198280
rect 148416 198228 148468 198280
rect 169024 198228 169076 198280
rect 169208 198228 169260 198280
rect 189172 198228 189224 198280
rect 106188 198092 106240 198144
rect 100576 198024 100628 198076
rect 61384 197956 61436 198008
rect 99288 197956 99340 198008
rect 127164 197956 127216 198008
rect 122196 197888 122248 197940
rect 131764 197888 131816 197940
rect 135996 198024 136048 198076
rect 142252 198092 142304 198144
rect 143448 198092 143500 198144
rect 164240 198160 164292 198212
rect 171784 198160 171836 198212
rect 172980 198160 173032 198212
rect 178408 198160 178460 198212
rect 208400 198160 208452 198212
rect 152924 198092 152976 198144
rect 154672 198092 154724 198144
rect 155960 198092 156012 198144
rect 162768 198024 162820 198076
rect 165436 198024 165488 198076
rect 169300 198092 169352 198144
rect 172244 198092 172296 198144
rect 173900 198092 173952 198144
rect 182180 198092 182232 198144
rect 219532 198092 219584 198144
rect 220728 198092 220780 198144
rect 169392 198024 169444 198076
rect 219440 198024 219492 198076
rect 138020 197956 138072 198008
rect 143448 197956 143500 198008
rect 146944 197956 146996 198008
rect 133972 197888 134024 197940
rect 139584 197888 139636 197940
rect 144184 197888 144236 197940
rect 561312 197956 561364 198008
rect 162952 197888 163004 197940
rect 177488 197888 177540 197940
rect 138756 197820 138808 197872
rect 145932 197820 145984 197872
rect 152096 197820 152148 197872
rect 154764 197820 154816 197872
rect 127808 197752 127860 197804
rect 138204 197752 138256 197804
rect 145564 197752 145616 197804
rect 148232 197752 148284 197804
rect 149060 197752 149112 197804
rect 113180 197684 113232 197736
rect 131028 197684 131080 197736
rect 141424 197684 141476 197736
rect 133144 197616 133196 197668
rect 142620 197616 142672 197668
rect 148048 197616 148100 197668
rect 150808 197616 150860 197668
rect 133972 197548 134024 197600
rect 144460 197548 144512 197600
rect 160284 197752 160336 197804
rect 169392 197752 169444 197804
rect 177580 197752 177632 197804
rect 178224 197752 178276 197804
rect 157156 197684 157208 197736
rect 164240 197684 164292 197736
rect 172520 197684 172572 197736
rect 172888 197684 172940 197736
rect 161848 197616 161900 197668
rect 170588 197616 170640 197668
rect 171416 197616 171468 197668
rect 177580 197616 177632 197668
rect 170772 197548 170824 197600
rect 138020 197480 138072 197532
rect 138756 197480 138808 197532
rect 140044 197480 140096 197532
rect 147864 197480 147916 197532
rect 151636 197480 151688 197532
rect 153936 197480 153988 197532
rect 154948 197480 155000 197532
rect 155408 197480 155460 197532
rect 160836 197480 160888 197532
rect 165620 197480 165672 197532
rect 146760 197412 146812 197464
rect 147312 197412 147364 197464
rect 149060 197412 149112 197464
rect 150348 197412 150400 197464
rect 164976 197412 165028 197464
rect 168012 197412 168064 197464
rect 139492 197344 139544 197396
rect 143816 197344 143868 197396
rect 146668 197344 146720 197396
rect 147128 197344 147180 197396
rect 147956 197344 148008 197396
rect 150716 197344 150768 197396
rect 168656 197344 168708 197396
rect 171508 197344 171560 197396
rect 172704 197344 172756 197396
rect 108396 197276 108448 197328
rect 170864 197276 170916 197328
rect 220728 197344 220780 197396
rect 580172 197344 580224 197396
rect 192300 197276 192352 197328
rect 193128 197276 193180 197328
rect 97356 197208 97408 197260
rect 161388 197208 161440 197260
rect 164056 197208 164108 197260
rect 111156 197140 111208 197192
rect 170772 197208 170824 197260
rect 171968 197208 172020 197260
rect 172336 197208 172388 197260
rect 173348 197208 173400 197260
rect 173900 197208 173952 197260
rect 189632 197208 189684 197260
rect 209872 197208 209924 197260
rect 169760 197140 169812 197192
rect 171416 197140 171468 197192
rect 171600 197140 171652 197192
rect 192576 197140 192628 197192
rect 112444 197072 112496 197124
rect 104256 197004 104308 197056
rect 107292 197004 107344 197056
rect 132408 197004 132460 197056
rect 135904 197004 135956 197056
rect 136364 197004 136416 197056
rect 136456 197004 136508 197056
rect 136640 197004 136692 197056
rect 146668 197072 146720 197124
rect 148140 197072 148192 197124
rect 149244 197072 149296 197124
rect 149704 197072 149756 197124
rect 149796 197072 149848 197124
rect 150348 197072 150400 197124
rect 161480 197072 161532 197124
rect 191932 197072 191984 197124
rect 193128 197072 193180 197124
rect 209964 197072 210016 197124
rect 118332 196936 118384 196988
rect 149520 196936 149572 196988
rect 153108 196936 153160 196988
rect 153844 196936 153896 196988
rect 158536 197004 158588 197056
rect 159640 197004 159692 197056
rect 166080 197004 166132 197056
rect 200212 197004 200264 197056
rect 156420 196936 156472 196988
rect 171876 196936 171928 196988
rect 171968 196936 172020 196988
rect 208492 196936 208544 196988
rect 104808 196868 104860 196920
rect 138572 196868 138624 196920
rect 144828 196868 144880 196920
rect 147036 196868 147088 196920
rect 148324 196868 148376 196920
rect 148508 196868 148560 196920
rect 157248 196868 157300 196920
rect 157524 196868 157576 196920
rect 117964 196732 118016 196784
rect 158168 196800 158220 196852
rect 158260 196800 158312 196852
rect 170312 196868 170364 196920
rect 170864 196868 170916 196920
rect 174084 196868 174136 196920
rect 212724 196868 212776 196920
rect 159364 196800 159416 196852
rect 163504 196800 163556 196852
rect 167920 196800 167972 196852
rect 169208 196800 169260 196852
rect 170772 196800 170824 196852
rect 173348 196800 173400 196852
rect 212632 196800 212684 196852
rect 138756 196732 138808 196784
rect 141056 196732 141108 196784
rect 143540 196732 143592 196784
rect 144460 196732 144512 196784
rect 146392 196732 146444 196784
rect 146852 196732 146904 196784
rect 148140 196732 148192 196784
rect 148784 196732 148836 196784
rect 154672 196732 154724 196784
rect 155592 196732 155644 196784
rect 155684 196732 155736 196784
rect 155868 196732 155920 196784
rect 156144 196732 156196 196784
rect 156788 196732 156840 196784
rect 157524 196732 157576 196784
rect 158352 196732 158404 196784
rect 158996 196732 159048 196784
rect 160008 196732 160060 196784
rect 163136 196732 163188 196784
rect 214656 196732 214708 196784
rect 96528 196664 96580 196716
rect 124404 196664 124456 196716
rect 136364 196664 136416 196716
rect 136640 196664 136692 196716
rect 139584 196664 139636 196716
rect 140688 196664 140740 196716
rect 141976 196664 142028 196716
rect 143172 196664 143224 196716
rect 143724 196664 143776 196716
rect 144276 196664 144328 196716
rect 146760 196664 146812 196716
rect 147588 196664 147640 196716
rect 147680 196664 147732 196716
rect 148876 196664 148928 196716
rect 149520 196664 149572 196716
rect 150072 196664 150124 196716
rect 150532 196664 150584 196716
rect 151452 196664 151504 196716
rect 152832 196664 152884 196716
rect 215300 196664 215352 196716
rect 3148 196596 3200 196648
rect 167276 196596 167328 196648
rect 169024 196596 169076 196648
rect 169760 196596 169812 196648
rect 170036 196596 170088 196648
rect 170496 196596 170548 196648
rect 173348 196596 173400 196648
rect 174084 196596 174136 196648
rect 174360 196596 174412 196648
rect 185400 196596 185452 196648
rect 207112 196596 207164 196648
rect 563704 196596 563756 196648
rect 121276 196528 121328 196580
rect 125416 196528 125468 196580
rect 142160 196528 142212 196580
rect 144736 196528 144788 196580
rect 145196 196528 145248 196580
rect 145840 196528 145892 196580
rect 154856 196528 154908 196580
rect 155776 196528 155828 196580
rect 159088 196528 159140 196580
rect 159548 196528 159600 196580
rect 160192 196528 160244 196580
rect 160376 196528 160428 196580
rect 163688 196528 163740 196580
rect 164148 196528 164200 196580
rect 168472 196528 168524 196580
rect 169484 196528 169536 196580
rect 170128 196528 170180 196580
rect 171968 196528 172020 196580
rect 131856 196460 131908 196512
rect 140780 196460 140832 196512
rect 143724 196460 143776 196512
rect 144644 196460 144696 196512
rect 150716 196460 150768 196512
rect 151360 196460 151412 196512
rect 155040 196460 155092 196512
rect 155592 196460 155644 196512
rect 156052 196460 156104 196512
rect 156880 196460 156932 196512
rect 157708 196460 157760 196512
rect 160836 196460 160888 196512
rect 164056 196460 164108 196512
rect 178684 196460 178736 196512
rect 116492 196392 116544 196444
rect 141608 196392 141660 196444
rect 142436 196392 142488 196444
rect 144920 196392 144972 196444
rect 145840 196392 145892 196444
rect 158076 196392 158128 196444
rect 158536 196392 158588 196444
rect 161664 196392 161716 196444
rect 162952 196392 163004 196444
rect 163964 196392 164016 196444
rect 164424 196392 164476 196444
rect 164700 196392 164752 196444
rect 165988 196392 166040 196444
rect 166816 196392 166868 196444
rect 168564 196392 168616 196444
rect 168932 196392 168984 196444
rect 171140 196392 171192 196444
rect 172060 196392 172112 196444
rect 176292 196392 176344 196444
rect 178408 196392 178460 196444
rect 167000 196324 167052 196376
rect 172888 196324 172940 196376
rect 131948 196256 132000 196308
rect 138940 196256 138992 196308
rect 140320 196256 140372 196308
rect 141608 196256 141660 196308
rect 156604 196256 156656 196308
rect 156972 196256 157024 196308
rect 159456 196256 159508 196308
rect 173164 196256 173216 196308
rect 158168 196188 158220 196240
rect 159732 196188 159784 196240
rect 161480 196188 161532 196240
rect 162676 196188 162728 196240
rect 168748 196188 168800 196240
rect 169576 196188 169628 196240
rect 137192 196052 137244 196104
rect 137468 196052 137520 196104
rect 120172 195984 120224 196036
rect 121460 195984 121512 196036
rect 134432 195916 134484 195968
rect 135168 195916 135220 195968
rect 138480 196120 138532 196172
rect 153384 196120 153436 196172
rect 166172 196120 166224 196172
rect 176200 196120 176252 196172
rect 138112 196052 138164 196104
rect 139952 196052 140004 196104
rect 142344 196052 142396 196104
rect 142804 196052 142856 196104
rect 153568 196052 153620 196104
rect 161664 196052 161716 196104
rect 162400 196052 162452 196104
rect 167000 196052 167052 196104
rect 167368 196052 167420 196104
rect 173900 196052 173952 196104
rect 174084 196052 174136 196104
rect 174176 196052 174228 196104
rect 174820 196052 174872 196104
rect 148324 195984 148376 196036
rect 148968 195984 149020 196036
rect 191196 195984 191248 196036
rect 215300 195984 215352 196036
rect 215576 195984 215628 196036
rect 580356 195984 580408 196036
rect 138480 195916 138532 195968
rect 139952 195916 140004 195968
rect 140412 195916 140464 195968
rect 149612 195916 149664 195968
rect 149888 195916 149940 195968
rect 156052 195916 156104 195968
rect 157064 195916 157116 195968
rect 160468 195916 160520 195968
rect 161296 195916 161348 195968
rect 163320 195916 163372 195968
rect 193220 195916 193272 195968
rect 197452 195916 197504 195968
rect 108304 195848 108356 195900
rect 171324 195848 171376 195900
rect 192944 195848 192996 195900
rect 108488 195780 108540 195832
rect 174452 195780 174504 195832
rect 176292 195780 176344 195832
rect 108672 195712 108724 195764
rect 170864 195712 170916 195764
rect 173900 195712 173952 195764
rect 198832 195712 198884 195764
rect 212816 195712 212868 195764
rect 213828 195712 213880 195764
rect 117780 195644 117832 195696
rect 147220 195644 147272 195696
rect 147772 195644 147824 195696
rect 148508 195644 148560 195696
rect 154212 195644 154264 195696
rect 154488 195644 154540 195696
rect 165436 195644 165488 195696
rect 170772 195644 170824 195696
rect 174360 195644 174412 195696
rect 175004 195644 175056 195696
rect 207296 195644 207348 195696
rect 122104 195576 122156 195628
rect 148232 195576 148284 195628
rect 166356 195576 166408 195628
rect 200304 195576 200356 195628
rect 117044 195508 117096 195560
rect 149336 195508 149388 195560
rect 110236 195440 110288 195492
rect 135536 195440 135588 195492
rect 137376 195440 137428 195492
rect 137652 195440 137704 195492
rect 139400 195440 139452 195492
rect 140412 195440 140464 195492
rect 100484 195372 100536 195424
rect 133236 195372 133288 195424
rect 144000 195372 144052 195424
rect 144184 195372 144236 195424
rect 109684 195304 109736 195356
rect 157248 195508 157300 195560
rect 165712 195508 165764 195560
rect 166540 195508 166592 195560
rect 168840 195508 168892 195560
rect 170496 195508 170548 195560
rect 173072 195508 173124 195560
rect 173532 195508 173584 195560
rect 179328 195508 179380 195560
rect 215300 195508 215352 195560
rect 152004 195440 152056 195492
rect 153016 195440 153068 195492
rect 4804 195236 4856 195288
rect 161756 195236 161808 195288
rect 164884 195372 164936 195424
rect 165160 195372 165212 195424
rect 165712 195372 165764 195424
rect 166448 195372 166500 195424
rect 178132 195440 178184 195492
rect 215484 195440 215536 195492
rect 169668 195372 169720 195424
rect 176292 195372 176344 195424
rect 208584 195372 208636 195424
rect 214380 195372 214432 195424
rect 323584 195372 323636 195424
rect 175464 195304 175516 195356
rect 212540 195304 212592 195356
rect 213828 195304 213880 195356
rect 574744 195304 574796 195356
rect 165160 195236 165212 195288
rect 165344 195236 165396 195288
rect 165896 195236 165948 195288
rect 166724 195236 166776 195288
rect 167368 195236 167420 195288
rect 168288 195236 168340 195288
rect 169944 195236 169996 195288
rect 209780 195236 209832 195288
rect 580816 195236 580868 195288
rect 108856 195168 108908 195220
rect 133328 195168 133380 195220
rect 137928 195168 137980 195220
rect 130752 195100 130804 195152
rect 139492 195100 139544 195152
rect 140964 195100 141016 195152
rect 141332 195100 141384 195152
rect 145380 195100 145432 195152
rect 178040 195168 178092 195220
rect 150992 195100 151044 195152
rect 152740 195100 152792 195152
rect 158628 195100 158680 195152
rect 182824 195100 182876 195152
rect 164608 195032 164660 195084
rect 165528 195032 165580 195084
rect 169668 195032 169720 195084
rect 180156 195032 180208 195084
rect 142528 194964 142580 195016
rect 169944 194964 169996 195016
rect 170680 194964 170732 195016
rect 173900 194964 173952 195016
rect 174636 194964 174688 195016
rect 105728 194896 105780 194948
rect 174360 194896 174412 194948
rect 141148 194828 141200 194880
rect 141700 194828 141752 194880
rect 141884 194828 141936 194880
rect 142528 194828 142580 194880
rect 165068 194828 165120 194880
rect 165436 194828 165488 194880
rect 169024 194828 169076 194880
rect 178776 194828 178828 194880
rect 128636 194760 128688 194812
rect 132040 194760 132092 194812
rect 166540 194760 166592 194812
rect 171876 194760 171928 194812
rect 133236 194692 133288 194744
rect 141240 194692 141292 194744
rect 130660 194624 130712 194676
rect 140044 194624 140096 194676
rect 202236 194624 202288 194676
rect 214012 194624 214064 194676
rect 214380 194624 214432 194676
rect 96344 194556 96396 194608
rect 103612 194556 103664 194608
rect 104624 194556 104676 194608
rect 178040 194556 178092 194608
rect 580264 194556 580316 194608
rect 104348 194488 104400 194540
rect 157432 194488 157484 194540
rect 163228 194488 163280 194540
rect 163872 194488 163924 194540
rect 190000 194488 190052 194540
rect 191840 194488 191892 194540
rect 107016 194420 107068 194472
rect 114376 194420 114428 194472
rect 164792 194420 164844 194472
rect 190920 194420 190972 194472
rect 202972 194420 203024 194472
rect 132224 194352 132276 194404
rect 133420 194352 133472 194404
rect 207020 194352 207072 194404
rect 103152 194284 103204 194336
rect 177120 194284 177172 194336
rect 195980 194284 196032 194336
rect 204444 194284 204496 194336
rect 94596 194216 94648 194268
rect 167000 194216 167052 194268
rect 170404 194216 170456 194268
rect 189632 194216 189684 194268
rect 190000 194216 190052 194268
rect 103060 194148 103112 194200
rect 176016 194148 176068 194200
rect 104624 194080 104676 194132
rect 114744 194080 114796 194132
rect 118056 194080 118108 194132
rect 121368 194080 121420 194132
rect 153200 194080 153252 194132
rect 190092 194148 190144 194200
rect 205640 194148 205692 194200
rect 200488 194080 200540 194132
rect 114376 194012 114428 194064
rect 146208 194012 146260 194064
rect 157616 194012 157668 194064
rect 174544 194012 174596 194064
rect 177120 194012 177172 194064
rect 177856 194012 177908 194064
rect 203064 194012 203116 194064
rect 102600 193944 102652 193996
rect 126980 193944 127032 193996
rect 149336 193944 149388 193996
rect 149980 193944 150032 193996
rect 157984 193944 158036 193996
rect 196624 193944 196676 193996
rect 198832 193944 198884 193996
rect 502984 193944 503036 193996
rect 94596 193876 94648 193928
rect 103520 193876 103572 193928
rect 104348 193876 104400 193928
rect 104624 193876 104676 193928
rect 137100 193876 137152 193928
rect 146208 193876 146260 193928
rect 151820 193876 151872 193928
rect 162584 193876 162636 193928
rect 195980 193876 196032 193928
rect 580632 193876 580684 193928
rect 3424 193808 3476 193860
rect 114100 193808 114152 193860
rect 146668 193808 146720 193860
rect 120356 193740 120408 193792
rect 142068 193740 142120 193792
rect 171508 193740 171560 193792
rect 188620 193740 188672 193792
rect 122012 193672 122064 193724
rect 135812 193672 135864 193724
rect 165620 193672 165672 193724
rect 185584 193672 185636 193724
rect 152464 193604 152516 193656
rect 328460 193604 328512 193656
rect 148508 193536 148560 193588
rect 579804 193536 579856 193588
rect 90456 193468 90508 193520
rect 164884 193468 164936 193520
rect 164976 193468 165028 193520
rect 165620 193468 165672 193520
rect 114928 193400 114980 193452
rect 147680 193400 147732 193452
rect 157800 193400 157852 193452
rect 158352 193400 158404 193452
rect 178040 193332 178092 193384
rect 178868 193332 178920 193384
rect 96620 193264 96672 193316
rect 118700 193264 118752 193316
rect 104164 193196 104216 193248
rect 112812 193196 112864 193248
rect 124956 193196 125008 193248
rect 132316 193196 132368 193248
rect 134524 193196 134576 193248
rect 170496 193196 170548 193248
rect 188712 193196 188764 193248
rect 142160 193128 142212 193180
rect 580448 193128 580500 193180
rect 138020 193060 138072 193112
rect 140044 193060 140096 193112
rect 142988 193060 143040 193112
rect 576400 193060 576452 193112
rect 132316 192992 132368 193044
rect 145748 192992 145800 193044
rect 577596 192992 577648 193044
rect 132960 192924 133012 192976
rect 201500 192924 201552 192976
rect 109868 192856 109920 192908
rect 163688 192856 163740 192908
rect 172244 192856 172296 192908
rect 108120 192788 108172 192840
rect 138204 192788 138256 192840
rect 147680 192788 147732 192840
rect 148692 192788 148744 192840
rect 189448 192788 189500 192840
rect 194692 192788 194744 192840
rect 204720 192788 204772 192840
rect 113088 192720 113140 192772
rect 146300 192720 146352 192772
rect 152188 192720 152240 192772
rect 152740 192720 152792 192772
rect 174268 192720 174320 192772
rect 208400 192720 208452 192772
rect 103336 192652 103388 192704
rect 135444 192652 135496 192704
rect 142436 192652 142488 192704
rect 332600 192652 332652 192704
rect 93308 192584 93360 192636
rect 101864 192584 101916 192636
rect 136364 192584 136416 192636
rect 171692 192584 171744 192636
rect 217140 192584 217192 192636
rect 561128 192584 561180 192636
rect 86224 192516 86276 192568
rect 99012 192516 99064 192568
rect 128636 192516 128688 192568
rect 132316 192516 132368 192568
rect 132960 192516 133012 192568
rect 160836 192516 160888 192568
rect 173256 192516 173308 192568
rect 175096 192516 175148 192568
rect 214288 192516 214340 192568
rect 580908 192516 580960 192568
rect 3424 192448 3476 192500
rect 124220 192448 124272 192500
rect 125508 192448 125560 192500
rect 127624 192448 127676 192500
rect 147220 192448 147272 192500
rect 156788 192448 156840 192500
rect 197360 192448 197412 192500
rect 208400 192448 208452 192500
rect 208952 192448 209004 192500
rect 577872 192448 577924 192500
rect 116400 192380 116452 192432
rect 139768 192380 139820 192432
rect 175188 192380 175240 192432
rect 189724 192380 189776 192432
rect 118700 192312 118752 192364
rect 144092 192312 144144 192364
rect 114744 192244 114796 192296
rect 144828 192244 144880 192296
rect 109408 192176 109460 192228
rect 140044 192176 140096 192228
rect 101772 191836 101824 191888
rect 105636 191836 105688 191888
rect 100208 191768 100260 191820
rect 111984 191768 112036 191820
rect 136916 191768 136968 191820
rect 137652 191768 137704 191820
rect 141516 191768 141568 191820
rect 144276 191768 144328 191820
rect 579160 191768 579212 191820
rect 103244 191700 103296 191752
rect 134432 191700 134484 191752
rect 137192 191700 137244 191752
rect 137928 191700 137980 191752
rect 139400 191700 139452 191752
rect 140688 191700 140740 191752
rect 256700 191700 256752 191752
rect 93124 191632 93176 191684
rect 165436 191632 165488 191684
rect 102692 191564 102744 191616
rect 172612 191564 172664 191616
rect 188804 191564 188856 191616
rect 97448 191496 97500 191548
rect 111156 191496 111208 191548
rect 117228 191496 117280 191548
rect 161940 191496 161992 191548
rect 162676 191496 162728 191548
rect 176108 191496 176160 191548
rect 200856 191496 200908 191548
rect 97264 191428 97316 191480
rect 108672 191428 108724 191480
rect 142252 191428 142304 191480
rect 159640 191428 159692 191480
rect 185676 191428 185728 191480
rect 100208 191360 100260 191412
rect 133880 191360 133932 191412
rect 135536 191360 135588 191412
rect 136548 191360 136600 191412
rect 137100 191360 137152 191412
rect 137744 191360 137796 191412
rect 155316 191360 155368 191412
rect 186412 191360 186464 191412
rect 100116 191292 100168 191344
rect 117228 191292 117280 191344
rect 154488 191292 154540 191344
rect 162676 191292 162728 191344
rect 196164 191292 196216 191344
rect 94688 191224 94740 191276
rect 111800 191224 111852 191276
rect 115296 191224 115348 191276
rect 150348 191224 150400 191276
rect 80060 191156 80112 191208
rect 118608 191156 118660 191208
rect 153292 191156 153344 191208
rect 99104 191088 99156 191140
rect 139400 191088 139452 191140
rect 109776 191020 109828 191072
rect 119436 191020 119488 191072
rect 149060 191020 149112 191072
rect 107108 190952 107160 191004
rect 115296 190952 115348 191004
rect 132684 190952 132736 191004
rect 132868 190952 132920 191004
rect 134064 190952 134116 191004
rect 134800 190952 134852 191004
rect 135720 190952 135772 191004
rect 136456 190952 136508 191004
rect 115848 190884 115900 190936
rect 132684 190816 132736 190868
rect 133420 190816 133472 190868
rect 137008 190816 137060 190868
rect 137560 190816 137612 190868
rect 152096 190884 152148 190936
rect 193956 191224 194008 191276
rect 167000 191156 167052 191208
rect 209136 191156 209188 191208
rect 159916 191088 159968 191140
rect 183468 191088 183520 191140
rect 578884 191088 578936 191140
rect 155408 191020 155460 191072
rect 155868 191020 155920 191072
rect 167276 190952 167328 191004
rect 167552 190952 167604 191004
rect 136916 190748 136968 190800
rect 137376 190748 137428 190800
rect 130476 190680 130528 190732
rect 141516 190680 141568 190732
rect 137192 190612 137244 190664
rect 137836 190612 137888 190664
rect 8944 190476 8996 190528
rect 100208 190476 100260 190528
rect 108580 190476 108632 190528
rect 113180 190476 113232 190528
rect 168840 190476 168892 190528
rect 199200 190476 199252 190528
rect 136640 190408 136692 190460
rect 137284 190408 137336 190460
rect 582748 190408 582800 190460
rect 133236 190340 133288 190392
rect 153108 190340 153160 190392
rect 577688 190340 577740 190392
rect 91744 190272 91796 190324
rect 170496 190272 170548 190324
rect 171784 190272 171836 190324
rect 191012 190272 191064 190324
rect 111800 190204 111852 190256
rect 112720 190204 112772 190256
rect 146852 190204 146904 190256
rect 169392 190204 169444 190256
rect 194876 190204 194928 190256
rect 113180 190136 113232 190188
rect 113732 190136 113784 190188
rect 146576 190136 146628 190188
rect 163504 190136 163556 190188
rect 193680 190136 193732 190188
rect 111984 190068 112036 190120
rect 145840 190068 145892 190120
rect 156696 190068 156748 190120
rect 190920 190068 190972 190120
rect 111524 190000 111576 190052
rect 136272 190000 136324 190052
rect 160652 190000 160704 190052
rect 195152 190000 195204 190052
rect 109776 189932 109828 189984
rect 133972 189932 134024 189984
rect 157524 189932 157576 189984
rect 192484 189932 192536 189984
rect 119528 189864 119580 189916
rect 150532 189864 150584 189916
rect 174176 189864 174228 189916
rect 209228 189864 209280 189916
rect 260840 189864 260892 189916
rect 119712 189796 119764 189848
rect 150992 189796 151044 189848
rect 157248 189796 157300 189848
rect 192300 189796 192352 189848
rect 194876 189796 194928 189848
rect 572260 189796 572312 189848
rect 107384 189728 107436 189780
rect 139492 189728 139544 189780
rect 156420 189728 156472 189780
rect 186136 189728 186188 189780
rect 579068 189728 579120 189780
rect 97356 189660 97408 189712
rect 104900 189660 104952 189712
rect 149520 189660 149572 189712
rect 170312 189660 170364 189712
rect 193220 189660 193272 189712
rect 111248 189592 111300 189644
rect 142804 189592 142856 189644
rect 169300 189592 169352 189644
rect 189080 189592 189132 189644
rect 170772 189524 170824 189576
rect 189356 189524 189408 189576
rect 105820 189184 105872 189236
rect 111984 189116 112036 189168
rect 112444 189116 112496 189168
rect 136640 189116 136692 189168
rect 3424 189048 3476 189100
rect 158628 189048 158680 189100
rect 206468 189048 206520 189100
rect 579620 189048 579672 189100
rect 110420 188980 110472 189032
rect 139860 188980 139912 189032
rect 144644 188980 144696 189032
rect 570604 188980 570656 189032
rect 100024 188844 100076 188896
rect 122932 188844 122984 188896
rect 123760 188844 123812 188896
rect 132132 188844 132184 188896
rect 143448 188912 143500 188964
rect 568028 188912 568080 188964
rect 149704 188844 149756 188896
rect 563796 188844 563848 188896
rect 94780 188776 94832 188828
rect 126796 188776 126848 188828
rect 143448 188776 143500 188828
rect 449164 188776 449216 188828
rect 94872 188708 94924 188760
rect 110512 188708 110564 188760
rect 116860 188708 116912 188760
rect 149704 188708 149756 188760
rect 150900 188708 150952 188760
rect 269764 188708 269816 188760
rect 98736 188640 98788 188692
rect 179420 188640 179472 188692
rect 205824 188640 205876 188692
rect 100300 188572 100352 188624
rect 177212 188572 177264 188624
rect 207388 188572 207440 188624
rect 153108 188504 153160 188556
rect 156880 188504 156932 188556
rect 171048 188504 171100 188556
rect 206008 188504 206060 188556
rect 206468 188504 206520 188556
rect 95884 188436 95936 188488
rect 154396 188436 154448 188488
rect 177764 188436 177816 188488
rect 215852 188436 215904 188488
rect 89168 188368 89220 188420
rect 153108 188368 153160 188420
rect 53840 188300 53892 188352
rect 107200 188300 107252 188352
rect 110512 188300 110564 188352
rect 111432 188300 111484 188352
rect 145196 188300 145248 188352
rect 149520 188300 149572 188352
rect 152740 188300 152792 188352
rect 163228 188368 163280 188420
rect 187056 188368 187108 188420
rect 241520 188368 241572 188420
rect 527180 188300 527232 188352
rect 123760 188232 123812 188284
rect 155592 188232 155644 188284
rect 102784 188096 102836 188148
rect 172888 188232 172940 188284
rect 203432 188232 203484 188284
rect 142804 187960 142856 188012
rect 150900 187960 150952 188012
rect 105636 187756 105688 187808
rect 110420 187756 110472 187808
rect 132040 187756 132092 187808
rect 143448 187756 143500 187808
rect 154396 187756 154448 187808
rect 155132 187756 155184 187808
rect 109592 187688 109644 187740
rect 144644 187688 144696 187740
rect 91836 187620 91888 187672
rect 171968 187620 172020 187672
rect 172244 187620 172296 187672
rect 199384 187620 199436 187672
rect 200304 187620 200356 187672
rect 569224 187620 569276 187672
rect 84844 187552 84896 187604
rect 107200 187484 107252 187536
rect 136180 187484 136232 187536
rect 166632 187552 166684 187604
rect 201132 187552 201184 187604
rect 163596 187484 163648 187536
rect 164148 187484 164200 187536
rect 168932 187484 168984 187536
rect 201776 187484 201828 187536
rect 126244 187416 126296 187468
rect 126796 187416 126848 187468
rect 151084 187416 151136 187468
rect 167460 187416 167512 187468
rect 201684 187416 201736 187468
rect 115112 187348 115164 187400
rect 147036 187348 147088 187400
rect 166080 187348 166132 187400
rect 200580 187348 200632 187400
rect 201408 187348 201460 187400
rect 108948 187280 109000 187332
rect 142344 187280 142396 187332
rect 163688 187280 163740 187332
rect 198004 187280 198056 187332
rect 111616 187212 111668 187264
rect 145104 187212 145156 187264
rect 158628 187212 158680 187264
rect 193864 187212 193916 187264
rect 108580 187144 108632 187196
rect 143356 187144 143408 187196
rect 165528 187144 165580 187196
rect 203156 187144 203208 187196
rect 112628 187076 112680 187128
rect 146760 187076 146812 187128
rect 173440 187076 173492 187128
rect 211804 187076 211856 187128
rect 100300 187008 100352 187060
rect 134984 187008 135036 187060
rect 135812 187008 135864 187060
rect 136180 187008 136232 187060
rect 158352 187008 158404 187060
rect 181996 187008 182048 187060
rect 278044 187008 278096 187060
rect 90548 186940 90600 186992
rect 158628 186940 158680 186992
rect 162216 186940 162268 186992
rect 196532 186940 196584 186992
rect 201408 186940 201460 186992
rect 572076 186940 572128 186992
rect 164148 186872 164200 186924
rect 176752 186872 176804 186924
rect 177672 186804 177724 186856
rect 210240 186872 210292 186924
rect 130844 186328 130896 186380
rect 144184 186328 144236 186380
rect 144828 186328 144880 186380
rect 158628 186328 158680 186380
rect 160008 186328 160060 186380
rect 102876 186260 102928 186312
rect 104348 186260 104400 186312
rect 112352 186260 112404 186312
rect 145656 186260 145708 186312
rect 569408 186260 569460 186312
rect 138020 186192 138072 186244
rect 558460 186192 558512 186244
rect 90364 186124 90416 186176
rect 121552 186124 121604 186176
rect 144828 186124 144880 186176
rect 512000 186124 512052 186176
rect 8300 186056 8352 186108
rect 168748 186056 168800 186108
rect 97816 185988 97868 186040
rect 189264 185988 189316 186040
rect 89260 185920 89312 185972
rect 178408 185920 178460 185972
rect 86408 185852 86460 185904
rect 161756 185852 161808 185904
rect 162676 185852 162728 185904
rect 203340 185920 203392 185972
rect 211712 185852 211764 185904
rect 93216 185784 93268 185836
rect 164700 185784 164752 185836
rect 170404 185784 170456 185836
rect 173808 185784 173860 185836
rect 207020 185784 207072 185836
rect 107660 185716 107712 185768
rect 169208 185716 169260 185768
rect 211252 185716 211304 185768
rect 212448 185716 212500 185768
rect 248420 185716 248472 185768
rect 104348 185648 104400 185700
rect 138296 185648 138348 185700
rect 150716 185648 150768 185700
rect 218428 185648 218480 185700
rect 306380 185648 306432 185700
rect 98828 185580 98880 185632
rect 138020 185580 138072 185632
rect 147588 185580 147640 185632
rect 215944 185580 215996 185632
rect 566740 185580 566792 185632
rect 106832 185512 106884 185564
rect 108488 185512 108540 185564
rect 140412 185512 140464 185564
rect 160560 185512 160612 185564
rect 211344 185512 211396 185564
rect 212448 185512 212500 185564
rect 121552 185444 121604 185496
rect 121920 185444 121972 185496
rect 161480 185444 161532 185496
rect 3424 185104 3476 185156
rect 7564 185104 7616 185156
rect 175648 184968 175700 185020
rect 210424 184968 210476 185020
rect 168748 184900 168800 184952
rect 210148 184900 210200 184952
rect 110328 184832 110380 184884
rect 143816 184832 143868 184884
rect 144736 184832 144788 184884
rect 581828 184832 581880 184884
rect 144828 184764 144880 184816
rect 572352 184764 572404 184816
rect 98920 184696 98972 184748
rect 167644 184696 167696 184748
rect 168196 184696 168248 184748
rect 173348 184696 173400 184748
rect 204536 184696 204588 184748
rect 95976 184628 96028 184680
rect 164608 184628 164660 184680
rect 165528 184628 165580 184680
rect 169944 184628 169996 184680
rect 203892 184628 203944 184680
rect 101496 184560 101548 184612
rect 168748 184560 168800 184612
rect 172244 184560 172296 184612
rect 205732 184560 205784 184612
rect 99932 184492 99984 184544
rect 158168 184492 158220 184544
rect 170036 184492 170088 184544
rect 204628 184492 204680 184544
rect 121092 184424 121144 184476
rect 154856 184424 154908 184476
rect 164884 184424 164936 184476
rect 199016 184424 199068 184476
rect 105912 184356 105964 184408
rect 139676 184356 139728 184408
rect 165436 184356 165488 184408
rect 199292 184356 199344 184408
rect 110052 184288 110104 184340
rect 143908 184288 143960 184340
rect 165528 184288 165580 184340
rect 206100 184288 206152 184340
rect 109684 184220 109736 184272
rect 143724 184220 143776 184272
rect 144828 184220 144880 184272
rect 159088 184220 159140 184272
rect 181904 184220 181956 184272
rect 436100 184220 436152 184272
rect 109500 184152 109552 184204
rect 144736 184152 144788 184204
rect 158260 184152 158312 184204
rect 216956 184152 217008 184204
rect 563888 184152 563940 184204
rect 104348 184084 104400 184136
rect 135904 184084 135956 184136
rect 160468 184084 160520 184136
rect 190552 184084 190604 184136
rect 108764 184016 108816 184068
rect 139584 184016 139636 184068
rect 176752 184016 176804 184068
rect 204812 184016 204864 184068
rect 106096 183948 106148 184000
rect 135536 183948 135588 184000
rect 168748 183948 168800 184000
rect 188896 183948 188948 184000
rect 109960 183880 110012 183932
rect 144552 183880 144604 183932
rect 80704 183472 80756 183524
rect 178224 183472 178276 183524
rect 178408 183472 178460 183524
rect 101404 183404 101456 183456
rect 178316 183404 178368 183456
rect 96160 183336 96212 183388
rect 141148 183336 141200 183388
rect 156236 183336 156288 183388
rect 202880 183336 202932 183388
rect 213000 183336 213052 183388
rect 178224 183268 178276 183320
rect 212908 183268 212960 183320
rect 178316 183200 178368 183252
rect 213092 183200 213144 183252
rect 165988 183132 166040 183184
rect 207204 183132 207256 183184
rect 164516 183064 164568 183116
rect 219624 183064 219676 183116
rect 159824 182996 159876 183048
rect 219808 182996 219860 183048
rect 313280 182996 313332 183048
rect 156328 182928 156380 182980
rect 216680 182928 216732 182980
rect 566832 182928 566884 182980
rect 158536 182860 158588 182912
rect 215760 182860 215812 182912
rect 582380 182860 582432 182912
rect 86316 182792 86368 182844
rect 125692 182792 125744 182844
rect 139216 182792 139268 182844
rect 153384 182792 153436 182844
rect 214840 182792 214892 182844
rect 583024 182792 583076 182844
rect 218244 182452 218296 182504
rect 218428 182452 218480 182504
rect 107108 182180 107160 182232
rect 187516 182180 187568 182232
rect 191932 182180 191984 182232
rect 193128 182180 193180 182232
rect 143448 182112 143500 182164
rect 150624 182112 150676 182164
rect 561220 182112 561272 182164
rect 162676 182044 162728 182096
rect 189448 182044 189500 182096
rect 193128 182044 193180 182096
rect 580172 182044 580224 182096
rect 142068 181976 142120 182028
rect 213920 181976 213972 182028
rect 171232 181908 171284 181960
rect 205916 181908 205968 181960
rect 176844 181840 176896 181892
rect 211620 181840 211672 181892
rect 152924 181772 152976 181824
rect 189264 181772 189316 181824
rect 106004 181704 106056 181756
rect 137100 181704 137152 181756
rect 156144 181704 156196 181756
rect 215668 181704 215720 181756
rect 233240 181704 233292 181756
rect 104256 181636 104308 181688
rect 137928 181636 137980 181688
rect 159180 181636 159232 181688
rect 180708 181636 180760 181688
rect 356060 181636 356112 181688
rect 103152 181568 103204 181620
rect 137560 181568 137612 181620
rect 152004 181568 152056 181620
rect 218520 181568 218572 181620
rect 562416 181568 562468 181620
rect 108396 181500 108448 181552
rect 142436 181500 142488 181552
rect 149428 181500 149480 181552
rect 217416 181500 217468 181552
rect 564072 181500 564124 181552
rect 94780 181432 94832 181484
rect 117964 181432 118016 181484
rect 126888 181432 126940 181484
rect 552756 181432 552808 181484
rect 174084 181364 174136 181416
rect 208768 181364 208820 181416
rect 175464 181296 175516 181348
rect 210332 181296 210384 181348
rect 3424 180820 3476 180872
rect 94780 180820 94832 180872
rect 103060 180820 103112 180872
rect 127808 180820 127860 180872
rect 563980 180752 564032 180804
rect 124036 180616 124088 180668
rect 556804 180684 556856 180736
rect 136180 180616 136232 180668
rect 558552 180616 558604 180668
rect 137008 180548 137060 180600
rect 558368 180548 558420 180600
rect 120724 180480 120776 180532
rect 455420 180480 455472 180532
rect 136916 180412 136968 180464
rect 362960 180412 363012 180464
rect 121000 180276 121052 180328
rect 136180 180276 136232 180328
rect 117964 180208 118016 180260
rect 149336 180208 149388 180260
rect 102968 180140 103020 180192
rect 137008 180140 137060 180192
rect 167368 180140 167420 180192
rect 208860 180140 208912 180192
rect 102876 180072 102928 180124
rect 136916 180072 136968 180124
rect 168656 180072 168708 180124
rect 219716 180072 219768 180124
rect 127716 179324 127768 179376
rect 581644 179324 581696 179376
rect 133788 179256 133840 179308
rect 578976 179256 579028 179308
rect 138756 179188 138808 179240
rect 558184 179188 558236 179240
rect 124772 179120 124824 179172
rect 139032 179120 139084 179172
rect 405740 179120 405792 179172
rect 124036 179052 124088 179104
rect 321560 179052 321612 179104
rect 170404 178848 170456 178900
rect 203248 178848 203300 178900
rect 167644 178780 167696 178832
rect 201868 178780 201920 178832
rect 105728 178712 105780 178764
rect 132868 178712 132920 178764
rect 133788 178712 133840 178764
rect 161664 178712 161716 178764
rect 210056 178712 210108 178764
rect 577780 178712 577832 178764
rect 105544 178644 105596 178696
rect 138756 178644 138808 178696
rect 164424 178644 164476 178696
rect 180616 178644 180668 178696
rect 560944 178644 560996 178696
rect 133788 177964 133840 178016
rect 555424 177964 555476 178016
rect 131120 177896 131172 177948
rect 132408 177896 132460 177948
rect 554044 177896 554096 177948
rect 191196 177828 191248 177880
rect 580172 177828 580224 177880
rect 136548 177760 136600 177812
rect 358820 177760 358872 177812
rect 101588 177420 101640 177472
rect 131120 177420 131172 177472
rect 98920 177352 98972 177404
rect 132776 177352 132828 177404
rect 133788 177352 133840 177404
rect 101496 177284 101548 177336
rect 136548 177284 136600 177336
rect 100116 176672 100168 176724
rect 122196 176672 122248 176724
rect 136456 176604 136508 176656
rect 552848 176604 552900 176656
rect 140780 176536 140832 176588
rect 141056 176536 141108 176588
rect 555516 176536 555568 176588
rect 395344 176468 395396 176520
rect 120908 175992 120960 176044
rect 140780 175992 140832 176044
rect 101680 175924 101732 175976
rect 136456 175924 136508 175976
rect 94872 173136 94924 173188
rect 116492 173136 116544 173188
rect 185676 173136 185728 173188
rect 580172 173136 580224 173188
rect 3424 172524 3476 172576
rect 94688 172524 94740 172576
rect 94872 172524 94924 172576
rect 116492 171776 116544 171828
rect 148784 171776 148836 171828
rect 110420 168988 110472 169040
rect 111156 168988 111208 169040
rect 116400 168988 116452 169040
rect 3148 168376 3200 168428
rect 110420 168376 110472 168428
rect 2780 165316 2832 165368
rect 4804 165316 4856 165368
rect 188344 164228 188396 164280
rect 580172 164228 580224 164280
rect 192576 162120 192628 162172
rect 206192 162120 206244 162172
rect 206192 161440 206244 161492
rect 580172 161440 580224 161492
rect 3516 161372 3568 161424
rect 171140 161372 171192 161424
rect 172244 161372 172296 161424
rect 172244 160692 172296 160744
rect 191932 160692 191984 160744
rect 3516 155932 3568 155984
rect 116952 155932 117004 155984
rect 127624 155864 127676 155916
rect 163136 153824 163188 153876
rect 198096 153824 198148 153876
rect 198096 153212 198148 153264
rect 579620 153212 579672 153264
rect 113548 153144 113600 153196
rect 117780 153144 117832 153196
rect 3516 151784 3568 151836
rect 113548 151784 113600 151836
rect 99932 151240 99984 151292
rect 132684 151240 132736 151292
rect 175464 151240 175516 151292
rect 210608 151240 210660 151292
rect 100024 151172 100076 151224
rect 134340 151172 134392 151224
rect 165896 151172 165948 151224
rect 217508 151172 217560 151224
rect 98644 151104 98696 151156
rect 132592 151104 132644 151156
rect 154764 151104 154816 151156
rect 214564 151104 214616 151156
rect 99840 151036 99892 151088
rect 134064 151036 134116 151088
rect 156052 151036 156104 151088
rect 216036 151036 216088 151088
rect 214656 149676 214708 149728
rect 580172 149676 580224 149728
rect 3424 148996 3476 149048
rect 160376 148996 160428 149048
rect 106924 148928 106976 148980
rect 132316 148928 132368 148980
rect 173992 148996 174044 149048
rect 207664 148996 207716 149048
rect 194784 148928 194836 148980
rect 106832 148860 106884 148912
rect 132224 148860 132276 148912
rect 165252 148860 165304 148912
rect 199660 148860 199712 148912
rect 104072 148792 104124 148844
rect 133236 148792 133288 148844
rect 163044 148792 163096 148844
rect 198280 148792 198332 148844
rect 110696 148724 110748 148776
rect 144460 148724 144512 148776
rect 167276 148724 167328 148776
rect 201960 148724 202012 148776
rect 101220 148656 101272 148708
rect 134248 148656 134300 148708
rect 161572 148656 161624 148708
rect 196900 148656 196952 148708
rect 98736 148588 98788 148640
rect 132960 148588 133012 148640
rect 168104 148588 168156 148640
rect 202052 148588 202104 148640
rect 108304 148520 108356 148572
rect 142620 148520 142672 148572
rect 168564 148520 168616 148572
rect 203616 148520 203668 148572
rect 101404 148452 101456 148504
rect 135720 148452 135772 148504
rect 169852 148452 169904 148504
rect 204996 148452 205048 148504
rect 107016 148384 107068 148436
rect 144000 148384 144052 148436
rect 175372 148384 175424 148436
rect 211988 148384 212040 148436
rect 97908 148316 97960 148368
rect 131764 148316 131816 148368
rect 174636 148316 174688 148368
rect 211896 148316 211948 148368
rect 120816 148248 120868 148300
rect 141700 148248 141752 148300
rect 167184 148248 167236 148300
rect 200672 148248 200724 148300
rect 110788 148180 110840 148232
rect 130752 148180 130804 148232
rect 172336 148180 172388 148232
rect 202144 148180 202196 148232
rect 114836 148112 114888 148164
rect 130660 148112 130712 148164
rect 180248 148112 180300 148164
rect 192760 148112 192812 148164
rect 171876 147296 171928 147348
rect 189816 147296 189868 147348
rect 176200 147228 176252 147280
rect 196072 147228 196124 147280
rect 168012 147160 168064 147212
rect 194048 147160 194100 147212
rect 165804 147092 165856 147144
rect 201408 147092 201460 147144
rect 112168 147024 112220 147076
rect 140320 147024 140372 147076
rect 165712 147024 165764 147076
rect 206376 147024 206428 147076
rect 101312 146956 101364 147008
rect 135628 146956 135680 147008
rect 168380 146956 168432 147008
rect 210516 146956 210568 147008
rect 102692 146888 102744 146940
rect 137468 146888 137520 146940
rect 580172 146888 580224 146940
rect 183284 146820 183336 146872
rect 183468 146820 183520 146872
rect 200948 146276 201000 146328
rect 201408 146276 201460 146328
rect 580448 146276 580500 146328
rect 116676 146208 116728 146260
rect 129372 146208 129424 146260
rect 179880 146208 179932 146260
rect 197912 146208 197964 146260
rect 115204 146140 115256 146192
rect 127072 146140 127124 146192
rect 177580 146140 177632 146192
rect 199752 146140 199804 146192
rect 113456 146072 113508 146124
rect 130384 146072 130436 146124
rect 173992 146072 174044 146124
rect 199108 146072 199160 146124
rect 112536 146004 112588 146056
rect 131764 146004 131816 146056
rect 172612 146004 172664 146056
rect 197820 146004 197872 146056
rect 114192 145936 114244 145988
rect 134248 145936 134300 145988
rect 162952 145936 163004 145988
rect 188344 145936 188396 145988
rect 111708 145868 111760 145920
rect 135260 145868 135312 145920
rect 169852 145868 169904 145920
rect 198740 145868 198792 145920
rect 112904 145800 112956 145852
rect 144092 145800 144144 145852
rect 167368 145800 167420 145852
rect 198924 145800 198976 145852
rect 119252 145732 119304 145784
rect 153752 145732 153804 145784
rect 160376 145732 160428 145784
rect 193588 145732 193640 145784
rect 118148 145664 118200 145716
rect 151912 145664 151964 145716
rect 164332 145664 164384 145716
rect 197636 145664 197688 145716
rect 119620 145596 119672 145648
rect 154488 145596 154540 145648
rect 162400 145596 162452 145648
rect 195244 145596 195296 145648
rect 117872 145528 117924 145580
rect 152372 145528 152424 145580
rect 162492 145528 162544 145580
rect 196808 145528 196860 145580
rect 112904 145460 112956 145512
rect 124220 145460 124272 145512
rect 177304 145460 177356 145512
rect 192392 145460 192444 145512
rect 116216 145392 116268 145444
rect 122932 145392 122984 145444
rect 181444 145392 181496 145444
rect 196256 145392 196308 145444
rect 113824 145324 113876 145376
rect 125232 145324 125284 145376
rect 184940 145324 184992 145376
rect 196440 145324 196492 145376
rect 120632 145256 120684 145308
rect 121368 145256 121420 145308
rect 188252 144984 188304 145036
rect 188896 144984 188948 145036
rect 3424 144916 3476 144968
rect 119068 144916 119120 144968
rect 119252 144916 119304 144968
rect 3516 144848 3568 144900
rect 113916 144848 113968 144900
rect 114192 144848 114244 144900
rect 121828 144848 121880 144900
rect 138664 144848 138716 144900
rect 176660 144848 176712 144900
rect 196348 144848 196400 144900
rect 197544 144848 197596 144900
rect 197728 144848 197780 144900
rect 580264 144848 580316 144900
rect 110972 144780 111024 144832
rect 130568 144780 130620 144832
rect 175280 144780 175332 144832
rect 199568 144780 199620 144832
rect 114468 144712 114520 144764
rect 140136 144712 140188 144764
rect 166908 144712 166960 144764
rect 196256 144712 196308 144764
rect 114284 144644 114336 144696
rect 141792 144644 141844 144696
rect 157340 144644 157392 144696
rect 189540 144644 189592 144696
rect 115572 144576 115624 144628
rect 142896 144576 142948 144628
rect 158168 144576 158220 144628
rect 190828 144576 190880 144628
rect 117688 144508 117740 144560
rect 149888 144508 149940 144560
rect 160284 144508 160336 144560
rect 195520 144508 195572 144560
rect 116400 144440 116452 144492
rect 148416 144440 148468 144492
rect 160192 144440 160244 144492
rect 194876 144440 194928 144492
rect 114744 144372 114796 144424
rect 148876 144372 148928 144424
rect 161296 144372 161348 144424
rect 195612 144372 195664 144424
rect 111340 144304 111392 144356
rect 145196 144304 145248 144356
rect 158076 144304 158128 144356
rect 194232 144304 194284 144356
rect 111708 144236 111760 144288
rect 146300 144236 146352 144288
rect 155868 144236 155920 144288
rect 191840 144236 191892 144288
rect 112996 144168 113048 144220
rect 137928 144168 137980 144220
rect 188160 144168 188212 144220
rect 196256 144168 196308 144220
rect 197084 144168 197136 144220
rect 207572 144168 207624 144220
rect 114192 144100 114244 144152
rect 126980 144100 127032 144152
rect 177488 144100 177540 144152
rect 198188 144100 198240 144152
rect 187608 144032 187660 144084
rect 197544 144032 197596 144084
rect 97816 143556 97868 143608
rect 111064 143488 111116 143540
rect 121552 143624 121604 143676
rect 191104 143624 191156 143676
rect 534080 143624 534132 143676
rect 118424 143556 118476 143608
rect 123668 143556 123720 143608
rect 492680 143556 492732 143608
rect 115480 143420 115532 143472
rect 121460 143488 121512 143540
rect 122196 143488 122248 143540
rect 122288 143488 122340 143540
rect 127624 143488 127676 143540
rect 172520 143488 172572 143540
rect 173716 143488 173768 143540
rect 133512 143420 133564 143472
rect 115204 143352 115256 143404
rect 119896 143352 119948 143404
rect 98000 143216 98052 143268
rect 97264 142944 97316 142996
rect 115204 142944 115256 142996
rect 82820 142808 82872 142860
rect 116308 143216 116360 143268
rect 116676 143216 116728 143268
rect 121552 143352 121604 143404
rect 127716 143352 127768 143404
rect 127808 143352 127860 143404
rect 138572 143352 138624 143404
rect 179328 143352 179380 143404
rect 187608 143352 187660 143404
rect 121368 143284 121420 143336
rect 139400 143284 139452 143336
rect 181352 143284 181404 143336
rect 192024 143284 192076 143336
rect 115664 143148 115716 143200
rect 120448 143148 120500 143200
rect 122288 143216 122340 143268
rect 126980 143216 127032 143268
rect 147680 143216 147732 143268
rect 177212 143216 177264 143268
rect 195060 143216 195112 143268
rect 140964 143148 141016 143200
rect 175188 143148 175240 143200
rect 197636 143148 197688 143200
rect 118516 143080 118568 143132
rect 145932 143080 145984 143132
rect 163872 143080 163924 143132
rect 193496 143080 193548 143132
rect 120632 143012 120684 143064
rect 143540 143012 143592 143064
rect 162308 143012 162360 143064
rect 194968 143012 195020 143064
rect 116584 142944 116636 142996
rect 119896 142944 119948 142996
rect 119988 142944 120040 142996
rect 150900 142944 150952 142996
rect 155684 142944 155736 142996
rect 157340 142944 157392 142996
rect 159824 142944 159876 142996
rect 193772 142944 193824 142996
rect 270500 142944 270552 142996
rect 116768 142876 116820 142928
rect 149244 142876 149296 142928
rect 168932 142876 168984 142928
rect 192208 142876 192260 142928
rect 192392 142876 192444 142928
rect 580264 142876 580316 142928
rect 119804 142808 119856 142860
rect 119896 142808 119948 142860
rect 120080 142808 120132 142860
rect 121368 142808 121420 142860
rect 122288 142808 122340 142860
rect 153384 142808 153436 142860
rect 166448 142808 166500 142860
rect 169760 142808 169812 142860
rect 171048 142808 171100 142860
rect 191104 142808 191156 142860
rect 192116 142808 192168 142860
rect 580724 142808 580776 142860
rect 116676 142740 116728 142792
rect 118240 142740 118292 142792
rect 131120 142740 131172 142792
rect 173716 142740 173768 142792
rect 179696 142740 179748 142792
rect 117136 142672 117188 142724
rect 128544 142672 128596 142724
rect 176384 142672 176436 142724
rect 178592 142672 178644 142724
rect 115756 142604 115808 142656
rect 126060 142604 126112 142656
rect 131120 142604 131172 142656
rect 426440 142604 426492 142656
rect 119804 142536 119856 142588
rect 122288 142536 122340 142588
rect 154488 142536 154540 142588
rect 514760 142536 514812 142588
rect 173716 142468 173768 142520
rect 179420 142468 179472 142520
rect 179696 142468 179748 142520
rect 207848 142468 207900 142520
rect 142896 142400 142948 142452
rect 188988 142400 189040 142452
rect 59360 142332 59412 142384
rect 177212 142332 177264 142384
rect 187608 142332 187660 142384
rect 220820 142332 220872 142384
rect 152372 142264 152424 142316
rect 365720 142264 365772 142316
rect 161388 142128 161440 142180
rect 114284 141992 114336 142044
rect 119896 142060 119948 142112
rect 151452 142060 151504 142112
rect 193312 142060 193364 142112
rect 146668 141992 146720 142044
rect 173256 141992 173308 142044
rect 192116 141992 192168 142044
rect 119988 141924 120040 141976
rect 151544 141924 151596 141976
rect 172428 141924 172480 141976
rect 193404 141924 193456 141976
rect 105452 141856 105504 141908
rect 138480 141856 138532 141908
rect 158352 141856 158404 141908
rect 190736 141856 190788 141908
rect 115572 141788 115624 141840
rect 148508 141788 148560 141840
rect 156512 141788 156564 141840
rect 190644 141788 190696 141840
rect 118148 141720 118200 141772
rect 152280 141720 152332 141772
rect 158628 141720 158680 141772
rect 193772 141720 193824 141772
rect 115020 141652 115072 141704
rect 149796 141652 149848 141704
rect 156972 141652 157024 141704
rect 191196 141652 191248 141704
rect 113824 141584 113876 141636
rect 148324 141584 148376 141636
rect 153108 141584 153160 141636
rect 191104 141584 191156 141636
rect 95976 141516 96028 141568
rect 139952 141516 140004 141568
rect 165160 141516 165212 141568
rect 206284 141516 206336 141568
rect 117872 141448 117924 141500
rect 178132 141448 178184 141500
rect 190644 141448 190696 141500
rect 395344 141448 395396 141500
rect 106740 141380 106792 141432
rect 172520 141380 172572 141432
rect 174820 141380 174872 141432
rect 190828 141380 190880 141432
rect 193312 141380 193364 141432
rect 518900 141380 518952 141432
rect 3516 141312 3568 141364
rect 8944 141312 8996 141364
rect 115664 141312 115716 141364
rect 145564 141312 145616 141364
rect 174544 141312 174596 141364
rect 190644 141312 190696 141364
rect 119620 140836 119672 140888
rect 119896 140836 119948 140888
rect 4804 140768 4856 140820
rect 158352 140768 158404 140820
rect 117136 140632 117188 140684
rect 147864 140700 147916 140752
rect 151912 140700 151964 140752
rect 152556 140700 152608 140752
rect 164332 140700 164384 140752
rect 164976 140700 165028 140752
rect 182824 140700 182876 140752
rect 192392 140700 192444 140752
rect 119252 140632 119304 140684
rect 123208 140632 123260 140684
rect 185952 140632 186004 140684
rect 190736 140632 190788 140684
rect 114008 140564 114060 140616
rect 124864 140564 124916 140616
rect 180156 140564 180208 140616
rect 196716 140564 196768 140616
rect 115848 140496 115900 140548
rect 132040 140496 132092 140548
rect 178684 140496 178736 140548
rect 195336 140496 195388 140548
rect 112536 140428 112588 140480
rect 131856 140428 131908 140480
rect 180064 140428 180116 140480
rect 199108 140428 199160 140480
rect 110880 140360 110932 140412
rect 131948 140360 132000 140412
rect 178776 140360 178828 140412
rect 197820 140360 197872 140412
rect 102784 140292 102836 140344
rect 133144 140292 133196 140344
rect 173164 140292 173216 140344
rect 193496 140292 193548 140344
rect 113916 140224 113968 140276
rect 145472 140224 145524 140276
rect 163780 140224 163832 140276
rect 186320 140224 186372 140276
rect 123484 140156 123536 140208
rect 149612 140156 149664 140208
rect 169944 140156 169996 140208
rect 204904 140156 204956 140208
rect 103980 140088 104032 140140
rect 137192 140088 137244 140140
rect 154672 140088 154724 140140
rect 214748 140088 214800 140140
rect 97172 140020 97224 140072
rect 138388 140020 138440 140072
rect 155776 140020 155828 140072
rect 189540 140020 189592 140072
rect 193588 140020 193640 140072
rect 335360 140020 335412 140072
rect 116676 139952 116728 140004
rect 123484 139952 123536 140004
rect 146668 139952 146720 140004
rect 146944 139952 146996 140004
rect 185584 139952 185636 140004
rect 190460 139952 190512 140004
rect 185860 139884 185912 139936
rect 193588 139884 193640 139936
rect 188344 139816 188396 139868
rect 188896 139816 188948 139868
rect 119804 139544 119856 139596
rect 124956 139544 125008 139596
rect 214748 139408 214800 139460
rect 580448 139408 580500 139460
rect 116768 138660 116820 138712
rect 129004 139272 129056 139324
rect 170588 139272 170640 139324
rect 188252 139272 188304 139324
rect 192760 138864 192812 138916
rect 202236 138864 202288 138916
rect 205088 138796 205140 138848
rect 196440 138728 196492 138780
rect 188988 138660 189040 138712
rect 580632 138660 580684 138712
rect 188988 137776 189040 137828
rect 197544 137776 197596 137828
rect 200856 137096 200908 137148
rect 203708 137096 203760 137148
rect 3424 136620 3476 136672
rect 105360 136620 105412 136672
rect 108120 136620 108172 136672
rect 203708 136620 203760 136672
rect 580172 136620 580224 136672
rect 118240 135872 118292 135924
rect 119988 135872 120040 135924
rect 196624 124856 196676 124908
rect 206468 124856 206520 124908
rect 206468 124176 206520 124228
rect 580172 124176 580224 124228
rect 3148 121388 3200 121440
rect 106740 121388 106792 121440
rect 3240 117240 3292 117292
rect 103980 117240 104032 117292
rect 210608 112412 210660 112464
rect 580172 112412 580224 112464
rect 3424 111800 3476 111852
rect 113640 111800 113692 111852
rect 3424 108944 3476 108996
rect 102140 108944 102192 108996
rect 102600 108944 102652 108996
rect 102140 108264 102192 108316
rect 112260 108264 112312 108316
rect 194048 105408 194100 105460
rect 202328 105408 202380 105460
rect 3424 103504 3476 103556
rect 119160 103504 119212 103556
rect 3424 96636 3476 96688
rect 117780 96636 117832 96688
rect 119344 95140 119396 95192
rect 120540 95140 120592 95192
rect 3148 93780 3200 93832
rect 115020 93780 115072 93832
rect 115020 92488 115072 92540
rect 119344 92488 119396 92540
rect 191288 91060 191340 91112
rect 198188 91060 198240 91112
rect 189724 85144 189776 85196
rect 189724 84872 189776 84924
rect 189172 84804 189224 84856
rect 189632 84804 189684 84856
rect 3424 84192 3476 84244
rect 98552 84192 98604 84244
rect 189172 82084 189224 82136
rect 206468 82084 206520 82136
rect 188620 81676 188672 81728
rect 188896 81676 188948 81728
rect 3424 81336 3476 81388
rect 108304 81336 108356 81388
rect 194232 81064 194284 81116
rect 108304 80860 108356 80912
rect 120080 80860 120132 80912
rect 120908 80860 120960 80912
rect 105636 80792 105688 80844
rect 113548 80724 113600 80776
rect 112352 80656 112404 80708
rect 117964 80588 118016 80640
rect 131764 80656 131816 80708
rect 131856 80656 131908 80708
rect 132040 80656 132092 80708
rect 123576 80452 123628 80504
rect 131764 80452 131816 80504
rect 119620 80384 119672 80436
rect 126244 80384 126296 80436
rect 119252 80316 119304 80368
rect 126336 80316 126388 80368
rect 128452 80316 128504 80368
rect 131856 80316 131908 80368
rect 128636 80248 128688 80300
rect 128544 80180 128596 80232
rect 132224 80180 132276 80232
rect 132040 80112 132092 80164
rect 124588 79976 124640 80028
rect 125232 79840 125284 79892
rect 132546 79908 132598 79960
rect 132914 79908 132966 79960
rect 133006 79908 133058 79960
rect 133374 79908 133426 79960
rect 133926 79908 133978 79960
rect 101220 79704 101272 79756
rect 97540 79636 97592 79688
rect 129004 79636 129056 79688
rect 132592 79704 132644 79756
rect 133282 79772 133334 79824
rect 115112 79568 115164 79620
rect 122840 79568 122892 79620
rect 131304 79568 131356 79620
rect 133144 79636 133196 79688
rect 133834 79840 133886 79892
rect 133558 79772 133610 79824
rect 133650 79772 133702 79824
rect 133512 79636 133564 79688
rect 133696 79636 133748 79688
rect 134110 79908 134162 79960
rect 134478 79908 134530 79960
rect 133972 79772 134024 79824
rect 113824 79500 113876 79552
rect 127532 79500 127584 79552
rect 96068 79432 96120 79484
rect 129280 79432 129332 79484
rect 121184 79364 121236 79416
rect 133328 79364 133380 79416
rect 133788 79364 133840 79416
rect 134294 79840 134346 79892
rect 135398 79908 135450 79960
rect 135490 79908 135542 79960
rect 135674 79908 135726 79960
rect 134202 79772 134254 79824
rect 134662 79772 134714 79824
rect 134846 79772 134898 79824
rect 135030 79772 135082 79824
rect 135214 79772 135266 79824
rect 134156 79636 134208 79688
rect 134432 79636 134484 79688
rect 135260 79636 135312 79688
rect 135352 79636 135404 79688
rect 134248 79432 134300 79484
rect 134984 79568 135036 79620
rect 134708 79500 134760 79552
rect 135950 79908 136002 79960
rect 136134 79908 136186 79960
rect 136226 79908 136278 79960
rect 136318 79908 136370 79960
rect 135904 79772 135956 79824
rect 136180 79704 136232 79756
rect 135628 79636 135680 79688
rect 135996 79636 136048 79688
rect 135904 79568 135956 79620
rect 136502 79908 136554 79960
rect 136870 79908 136922 79960
rect 137054 79908 137106 79960
rect 136456 79636 136508 79688
rect 137146 79840 137198 79892
rect 137100 79704 137152 79756
rect 136364 79568 136416 79620
rect 136916 79568 136968 79620
rect 137008 79568 137060 79620
rect 137606 79908 137658 79960
rect 137790 79908 137842 79960
rect 137882 79908 137934 79960
rect 138066 79908 138118 79960
rect 138158 79908 138210 79960
rect 137468 79568 137520 79620
rect 138342 79840 138394 79892
rect 138526 79840 138578 79892
rect 138112 79772 138164 79824
rect 138710 79908 138762 79960
rect 138986 79908 139038 79960
rect 138802 79840 138854 79892
rect 138894 79840 138946 79892
rect 139078 79772 139130 79824
rect 138756 79704 138808 79756
rect 138940 79704 138992 79756
rect 138572 79636 138624 79688
rect 139032 79636 139084 79688
rect 137836 79568 137888 79620
rect 137928 79568 137980 79620
rect 138020 79568 138072 79620
rect 138848 79568 138900 79620
rect 139538 79908 139590 79960
rect 139906 79908 139958 79960
rect 139998 79908 140050 79960
rect 141102 79908 141154 79960
rect 140550 79840 140602 79892
rect 140826 79840 140878 79892
rect 140044 79772 140096 79824
rect 139492 79704 139544 79756
rect 141194 79840 141246 79892
rect 141286 79840 141338 79892
rect 141654 79908 141706 79960
rect 141930 79908 141982 79960
rect 142114 79908 142166 79960
rect 142390 79908 142442 79960
rect 142482 79908 142534 79960
rect 141838 79840 141890 79892
rect 141148 79704 141200 79756
rect 141470 79772 141522 79824
rect 141562 79772 141614 79824
rect 139400 79636 139452 79688
rect 140780 79636 140832 79688
rect 141056 79636 141108 79688
rect 141332 79636 141384 79688
rect 141424 79636 141476 79688
rect 141516 79636 141568 79688
rect 141608 79636 141660 79688
rect 141884 79704 141936 79756
rect 140412 79568 140464 79620
rect 142758 79840 142810 79892
rect 142574 79772 142626 79824
rect 142436 79636 142488 79688
rect 142528 79636 142580 79688
rect 142620 79636 142672 79688
rect 142252 79568 142304 79620
rect 143126 79908 143178 79960
rect 143402 79908 143454 79960
rect 143080 79636 143132 79688
rect 143356 79568 143408 79620
rect 144138 79908 144190 79960
rect 144230 79908 144282 79960
rect 144322 79908 144374 79960
rect 143678 79840 143730 79892
rect 143770 79840 143822 79892
rect 143954 79840 144006 79892
rect 144046 79840 144098 79892
rect 143632 79636 143684 79688
rect 143908 79568 143960 79620
rect 144184 79704 144236 79756
rect 144184 79568 144236 79620
rect 144506 79840 144558 79892
rect 144598 79840 144650 79892
rect 144460 79636 144512 79688
rect 144552 79568 144604 79620
rect 188620 80996 188672 81048
rect 202880 80996 202932 81048
rect 203708 80928 203760 80980
rect 207388 80860 207440 80912
rect 177856 80656 177908 80708
rect 177948 80656 178000 80708
rect 195336 80724 195388 80776
rect 182824 80656 182876 80708
rect 211988 80656 212040 80708
rect 144874 79908 144926 79960
rect 144966 79908 145018 79960
rect 145058 79908 145110 79960
rect 145150 79908 145202 79960
rect 145426 79908 145478 79960
rect 145794 79908 145846 79960
rect 145978 79908 146030 79960
rect 146070 79908 146122 79960
rect 146438 79908 146490 79960
rect 146622 79908 146674 79960
rect 146898 79908 146950 79960
rect 147266 79908 147318 79960
rect 147358 79908 147410 79960
rect 144828 79772 144880 79824
rect 145104 79772 145156 79824
rect 145196 79772 145248 79824
rect 144920 79704 144972 79756
rect 145012 79636 145064 79688
rect 145702 79840 145754 79892
rect 145656 79704 145708 79756
rect 145748 79704 145800 79756
rect 145932 79704 145984 79756
rect 146254 79840 146306 79892
rect 146116 79704 146168 79756
rect 146208 79704 146260 79756
rect 146392 79704 146444 79756
rect 146024 79636 146076 79688
rect 146806 79840 146858 79892
rect 145564 79568 145616 79620
rect 136732 79500 136784 79552
rect 134892 79432 134944 79484
rect 140780 79432 140832 79484
rect 142804 79500 142856 79552
rect 143540 79500 143592 79552
rect 143816 79500 143868 79552
rect 144092 79500 144144 79552
rect 145472 79500 145524 79552
rect 145840 79500 145892 79552
rect 146668 79500 146720 79552
rect 147312 79772 147364 79824
rect 147542 79908 147594 79960
rect 147726 79908 147778 79960
rect 148462 79908 148514 79960
rect 148738 79908 148790 79960
rect 148922 79908 148974 79960
rect 149198 79908 149250 79960
rect 149382 79908 149434 79960
rect 149658 79908 149710 79960
rect 149842 79908 149894 79960
rect 149934 79908 149986 79960
rect 150486 79908 150538 79960
rect 147404 79704 147456 79756
rect 147910 79840 147962 79892
rect 148094 79840 148146 79892
rect 148186 79840 148238 79892
rect 147680 79772 147732 79824
rect 146944 79636 146996 79688
rect 147496 79636 147548 79688
rect 147956 79568 148008 79620
rect 148370 79772 148422 79824
rect 148232 79636 148284 79688
rect 148508 79636 148560 79688
rect 148600 79636 148652 79688
rect 148830 79840 148882 79892
rect 148876 79636 148928 79688
rect 149566 79840 149618 79892
rect 148232 79500 148284 79552
rect 149060 79568 149112 79620
rect 148968 79500 149020 79552
rect 149428 79636 149480 79688
rect 149244 79568 149296 79620
rect 149612 79636 149664 79688
rect 149796 79568 149848 79620
rect 150302 79840 150354 79892
rect 150256 79704 150308 79756
rect 150440 79704 150492 79756
rect 149704 79500 149756 79552
rect 151038 79908 151090 79960
rect 151130 79908 151182 79960
rect 151314 79908 151366 79960
rect 151406 79908 151458 79960
rect 151590 79908 151642 79960
rect 150762 79840 150814 79892
rect 151268 79772 151320 79824
rect 151544 79636 151596 79688
rect 150808 79568 150860 79620
rect 151084 79568 151136 79620
rect 188344 80588 188396 80640
rect 189908 80588 189960 80640
rect 152418 79908 152470 79960
rect 152786 79908 152838 79960
rect 152878 79908 152930 79960
rect 153154 79908 153206 79960
rect 153430 79908 153482 79960
rect 154166 79908 154218 79960
rect 154258 79908 154310 79960
rect 154626 79908 154678 79960
rect 154902 79908 154954 79960
rect 154994 79908 155046 79960
rect 155086 79908 155138 79960
rect 155270 79908 155322 79960
rect 155362 79908 155414 79960
rect 155638 79908 155690 79960
rect 155730 79908 155782 79960
rect 155822 79908 155874 79960
rect 155914 79908 155966 79960
rect 156006 79908 156058 79960
rect 156098 79908 156150 79960
rect 156190 79908 156242 79960
rect 156374 79908 156426 79960
rect 156650 79908 156702 79960
rect 156926 79908 156978 79960
rect 157202 79908 157254 79960
rect 157294 79908 157346 79960
rect 158122 79908 158174 79960
rect 158490 79908 158542 79960
rect 158582 79908 158634 79960
rect 158674 79908 158726 79960
rect 159318 79908 159370 79960
rect 159410 79908 159462 79960
rect 159686 79908 159738 79960
rect 159870 79908 159922 79960
rect 159962 79908 160014 79960
rect 160054 79908 160106 79960
rect 151958 79840 152010 79892
rect 152050 79840 152102 79892
rect 152234 79840 152286 79892
rect 150716 79500 150768 79552
rect 151636 79500 151688 79552
rect 151820 79500 151872 79552
rect 3516 79296 3568 79348
rect 140780 79296 140832 79348
rect 112260 79228 112312 79280
rect 134432 79228 134484 79280
rect 139492 79228 139544 79280
rect 140504 79228 140556 79280
rect 141424 79364 141476 79416
rect 151176 79364 151228 79416
rect 151912 79364 151964 79416
rect 152188 79704 152240 79756
rect 152694 79840 152746 79892
rect 152648 79704 152700 79756
rect 152970 79840 153022 79892
rect 153016 79704 153068 79756
rect 153246 79840 153298 79892
rect 152648 79432 152700 79484
rect 152832 79636 152884 79688
rect 152924 79636 152976 79688
rect 153108 79636 153160 79688
rect 153798 79840 153850 79892
rect 153982 79840 154034 79892
rect 153476 79704 153528 79756
rect 153936 79704 153988 79756
rect 153384 79636 153436 79688
rect 153752 79636 153804 79688
rect 154120 79704 154172 79756
rect 154810 79840 154862 79892
rect 154856 79704 154908 79756
rect 154580 79636 154632 79688
rect 154764 79636 154816 79688
rect 154672 79568 154724 79620
rect 153936 79432 153988 79484
rect 154304 79364 154356 79416
rect 155132 79636 155184 79688
rect 155454 79772 155506 79824
rect 155592 79772 155644 79824
rect 155914 79772 155966 79824
rect 155776 79704 155828 79756
rect 155500 79636 155552 79688
rect 155684 79636 155736 79688
rect 155868 79636 155920 79688
rect 156144 79704 156196 79756
rect 155408 79568 155460 79620
rect 156466 79772 156518 79824
rect 156328 79636 156380 79688
rect 156512 79636 156564 79688
rect 156420 79568 156472 79620
rect 155960 79500 156012 79552
rect 156604 79500 156656 79552
rect 157478 79840 157530 79892
rect 157938 79840 157990 79892
rect 157248 79704 157300 79756
rect 157616 79704 157668 79756
rect 158168 79772 158220 79824
rect 157984 79636 158036 79688
rect 157616 79568 157668 79620
rect 157708 79500 157760 79552
rect 157340 79432 157392 79484
rect 141240 79296 141292 79348
rect 152464 79296 152516 79348
rect 157432 79296 157484 79348
rect 158444 79568 158496 79620
rect 158766 79772 158818 79824
rect 158812 79636 158864 79688
rect 159364 79704 159416 79756
rect 158536 79500 158588 79552
rect 158260 79432 158312 79484
rect 158904 79500 158956 79552
rect 158996 79500 159048 79552
rect 158904 79364 158956 79416
rect 159594 79772 159646 79824
rect 159548 79636 159600 79688
rect 159640 79568 159692 79620
rect 160330 79908 160382 79960
rect 160422 79908 160474 79960
rect 160514 79908 160566 79960
rect 160606 79908 160658 79960
rect 160698 79908 160750 79960
rect 160790 79908 160842 79960
rect 160882 79908 160934 79960
rect 161066 79908 161118 79960
rect 161434 79908 161486 79960
rect 161618 79908 161670 79960
rect 161710 79908 161762 79960
rect 161802 79908 161854 79960
rect 161986 79908 162038 79960
rect 162446 79908 162498 79960
rect 162538 79908 162590 79960
rect 162814 79908 162866 79960
rect 162998 79908 163050 79960
rect 163090 79908 163142 79960
rect 163274 79908 163326 79960
rect 160192 79568 160244 79620
rect 159824 79500 159876 79552
rect 160008 79500 160060 79552
rect 160514 79772 160566 79824
rect 160468 79636 160520 79688
rect 161112 79704 161164 79756
rect 160836 79636 160888 79688
rect 161894 79840 161946 79892
rect 161756 79704 161808 79756
rect 161848 79704 161900 79756
rect 160652 79568 160704 79620
rect 161204 79568 161256 79620
rect 161664 79568 161716 79620
rect 161572 79500 161624 79552
rect 162492 79704 162544 79756
rect 162722 79772 162774 79824
rect 162676 79636 162728 79688
rect 162768 79568 162820 79620
rect 162032 79500 162084 79552
rect 163044 79772 163096 79824
rect 163642 79908 163694 79960
rect 163826 79908 163878 79960
rect 164102 79908 164154 79960
rect 164562 79908 164614 79960
rect 164654 79908 164706 79960
rect 164746 79908 164798 79960
rect 164930 79908 164982 79960
rect 165022 79908 165074 79960
rect 165206 79908 165258 79960
rect 165390 79908 165442 79960
rect 165666 79908 165718 79960
rect 165758 79908 165810 79960
rect 163412 79636 163464 79688
rect 163734 79840 163786 79892
rect 163872 79772 163924 79824
rect 164378 79840 164430 79892
rect 164194 79772 164246 79824
rect 163688 79636 163740 79688
rect 164056 79636 164108 79688
rect 164240 79636 164292 79688
rect 164516 79704 164568 79756
rect 163596 79568 163648 79620
rect 164424 79568 164476 79620
rect 164608 79568 164660 79620
rect 165344 79772 165396 79824
rect 164976 79704 165028 79756
rect 165160 79704 165212 79756
rect 164884 79636 164936 79688
rect 165574 79840 165626 79892
rect 165620 79704 165672 79756
rect 165942 79840 165994 79892
rect 165804 79704 165856 79756
rect 166126 79772 166178 79824
rect 165896 79636 165948 79688
rect 166080 79636 166132 79688
rect 165436 79568 165488 79620
rect 166402 79908 166454 79960
rect 166494 79908 166546 79960
rect 166678 79908 166730 79960
rect 166770 79908 166822 79960
rect 167138 79908 167190 79960
rect 167230 79908 167282 79960
rect 167506 79908 167558 79960
rect 167690 79908 167742 79960
rect 167782 79908 167834 79960
rect 168426 79908 168478 79960
rect 168794 79908 168846 79960
rect 168886 79908 168938 79960
rect 168978 79908 169030 79960
rect 169070 79908 169122 79960
rect 169346 79908 169398 79960
rect 166310 79772 166362 79824
rect 166632 79704 166684 79756
rect 166356 79636 166408 79688
rect 166448 79636 166500 79688
rect 166540 79568 166592 79620
rect 167322 79840 167374 79892
rect 167276 79704 167328 79756
rect 167598 79840 167650 79892
rect 167460 79636 167512 79688
rect 167000 79568 167052 79620
rect 167184 79568 167236 79620
rect 167368 79568 167420 79620
rect 167552 79568 167604 79620
rect 163320 79500 163372 79552
rect 164700 79500 164752 79552
rect 168518 79840 168570 79892
rect 168472 79636 168524 79688
rect 168932 79772 168984 79824
rect 168840 79704 168892 79756
rect 167828 79568 167880 79620
rect 168564 79568 168616 79620
rect 169024 79568 169076 79620
rect 186964 80520 187016 80572
rect 192668 80520 192720 80572
rect 179604 80452 179656 80504
rect 187056 80452 187108 80504
rect 191104 80452 191156 80504
rect 178132 80384 178184 80436
rect 178040 80248 178092 80300
rect 169714 79908 169766 79960
rect 169898 79908 169950 79960
rect 170174 79908 170226 79960
rect 170450 79908 170502 79960
rect 170542 79908 170594 79960
rect 171278 79908 171330 79960
rect 171646 79908 171698 79960
rect 172106 79908 172158 79960
rect 172198 79908 172250 79960
rect 172382 79908 172434 79960
rect 172566 79908 172618 79960
rect 173026 79908 173078 79960
rect 169668 79772 169720 79824
rect 170358 79840 170410 79892
rect 170312 79704 170364 79756
rect 170404 79704 170456 79756
rect 171002 79840 171054 79892
rect 171186 79840 171238 79892
rect 170036 79636 170088 79688
rect 170128 79636 170180 79688
rect 170496 79636 170548 79688
rect 170956 79636 171008 79688
rect 169392 79568 169444 79620
rect 167920 79500 167972 79552
rect 165620 79432 165672 79484
rect 162584 79364 162636 79416
rect 141424 79228 141476 79280
rect 145288 79228 145340 79280
rect 145564 79228 145616 79280
rect 166540 79364 166592 79416
rect 168288 79364 168340 79416
rect 171830 79840 171882 79892
rect 171600 79636 171652 79688
rect 171968 79636 172020 79688
rect 177764 80180 177816 80232
rect 178960 80180 179012 80232
rect 179236 80044 179288 80096
rect 203800 80044 203852 80096
rect 204720 80044 204772 80096
rect 182824 79976 182876 80028
rect 183928 79976 183980 80028
rect 190828 79976 190880 80028
rect 202328 79976 202380 80028
rect 202788 79976 202840 80028
rect 580172 79976 580224 80028
rect 173762 79908 173814 79960
rect 172428 79772 172480 79824
rect 172612 79772 172664 79824
rect 172244 79704 172296 79756
rect 172336 79636 172388 79688
rect 171784 79568 171836 79620
rect 173210 79840 173262 79892
rect 173578 79840 173630 79892
rect 173394 79772 173446 79824
rect 173440 79636 173492 79688
rect 174866 79908 174918 79960
rect 174958 79908 175010 79960
rect 175418 79908 175470 79960
rect 175878 79908 175930 79960
rect 174038 79840 174090 79892
rect 174130 79840 174182 79892
rect 173900 79636 173952 79688
rect 174498 79772 174550 79824
rect 174590 79772 174642 79824
rect 174912 79772 174964 79824
rect 174820 79636 174872 79688
rect 173256 79568 173308 79620
rect 173532 79568 173584 79620
rect 173624 79568 173676 79620
rect 173992 79568 174044 79620
rect 174544 79568 174596 79620
rect 175142 79840 175194 79892
rect 175326 79840 175378 79892
rect 175786 79840 175838 79892
rect 175510 79772 175562 79824
rect 175602 79772 175654 79824
rect 175372 79704 175424 79756
rect 175004 79636 175056 79688
rect 175280 79636 175332 79688
rect 175464 79636 175516 79688
rect 175832 79704 175884 79756
rect 176154 79908 176206 79960
rect 176246 79908 176298 79960
rect 176430 79908 176482 79960
rect 177856 79908 177908 79960
rect 185584 79908 185636 79960
rect 214288 79908 214340 79960
rect 176706 79840 176758 79892
rect 176798 79840 176850 79892
rect 176982 79840 177034 79892
rect 177074 79840 177126 79892
rect 177166 79840 177218 79892
rect 177764 79840 177816 79892
rect 176200 79772 176252 79824
rect 175648 79636 175700 79688
rect 176016 79636 176068 79688
rect 176292 79568 176344 79620
rect 171416 79364 171468 79416
rect 175924 79500 175976 79552
rect 176660 79568 176712 79620
rect 179052 79840 179104 79892
rect 178040 79704 178092 79756
rect 580632 79704 580684 79756
rect 177120 79568 177172 79620
rect 179788 79568 179840 79620
rect 176844 79500 176896 79552
rect 177028 79500 177080 79552
rect 177396 79500 177448 79552
rect 209136 79500 209188 79552
rect 172060 79432 172112 79484
rect 172704 79432 172756 79484
rect 173532 79432 173584 79484
rect 189172 79432 189224 79484
rect 119436 79160 119488 79212
rect 150348 79160 150400 79212
rect 112444 79092 112496 79144
rect 144920 79092 144972 79144
rect 145288 79092 145340 79144
rect 145748 79092 145800 79144
rect 151176 79092 151228 79144
rect 168104 79228 168156 79280
rect 201868 79364 201920 79416
rect 161480 79160 161532 79212
rect 170680 79160 170732 79212
rect 171048 79160 171100 79212
rect 173532 79296 173584 79348
rect 198004 79296 198056 79348
rect 118056 79024 118108 79076
rect 153016 79024 153068 79076
rect 111248 78956 111300 79008
rect 146116 78956 146168 79008
rect 149060 78956 149112 79008
rect 164240 79024 164292 79076
rect 172152 79160 172204 79212
rect 175372 79228 175424 79280
rect 175556 79228 175608 79280
rect 176292 79228 176344 79280
rect 176476 79228 176528 79280
rect 210424 79228 210476 79280
rect 174912 79160 174964 79212
rect 209228 79160 209280 79212
rect 181352 79092 181404 79144
rect 172888 78956 172940 79008
rect 174084 78956 174136 79008
rect 121920 78888 121972 78940
rect 162676 78888 162728 78940
rect 167920 78888 167972 78940
rect 181444 79024 181496 79076
rect 176752 78956 176804 79008
rect 210608 79092 210660 79144
rect 181628 78956 181680 79008
rect 202788 79024 202840 79076
rect 178132 78888 178184 78940
rect 212724 78888 212776 78940
rect 98828 78820 98880 78872
rect 139584 78820 139636 78872
rect 142344 78820 142396 78872
rect 142988 78820 143040 78872
rect 158352 78820 158404 78872
rect 158720 78820 158772 78872
rect 171140 78820 171192 78872
rect 211528 78820 211580 78872
rect 133328 78752 133380 78804
rect 137008 78752 137060 78804
rect 140504 78752 140556 78804
rect 144644 78752 144696 78804
rect 146116 78752 146168 78804
rect 148508 78752 148560 78804
rect 172336 78752 172388 78804
rect 217140 78752 217192 78804
rect 129648 78684 129700 78736
rect 138020 78684 138072 78736
rect 168380 78684 168432 78736
rect 172060 78684 172112 78736
rect 181352 78684 181404 78736
rect 182180 78684 182232 78736
rect 121000 78616 121052 78668
rect 135812 78616 135864 78668
rect 136640 78616 136692 78668
rect 143264 78616 143316 78668
rect 154580 78616 154632 78668
rect 154948 78616 155000 78668
rect 155592 78616 155644 78668
rect 158352 78616 158404 78668
rect 160100 78616 160152 78668
rect 160284 78616 160336 78668
rect 168656 78616 168708 78668
rect 169300 78616 169352 78668
rect 174084 78616 174136 78668
rect 188804 78616 188856 78668
rect 131028 78548 131080 78600
rect 138388 78548 138440 78600
rect 142620 78548 142672 78600
rect 142804 78548 142856 78600
rect 167000 78548 167052 78600
rect 168196 78548 168248 78600
rect 173072 78548 173124 78600
rect 209964 78548 210016 78600
rect 104532 78480 104584 78532
rect 127440 78480 127492 78532
rect 131856 78480 131908 78532
rect 141516 78480 141568 78532
rect 175924 78480 175976 78532
rect 207848 78480 207900 78532
rect 104072 78412 104124 78464
rect 129648 78412 129700 78464
rect 131120 78412 131172 78464
rect 132316 78412 132368 78464
rect 132500 78412 132552 78464
rect 136732 78412 136784 78464
rect 155868 78412 155920 78464
rect 156604 78412 156656 78464
rect 166540 78412 166592 78464
rect 104440 78344 104492 78396
rect 128544 78344 128596 78396
rect 131212 78344 131264 78396
rect 138940 78344 138992 78396
rect 140412 78344 140464 78396
rect 147404 78344 147456 78396
rect 163228 78344 163280 78396
rect 166632 78344 166684 78396
rect 171784 78412 171836 78464
rect 206192 78412 206244 78464
rect 188896 78344 188948 78396
rect 106832 78276 106884 78328
rect 131304 78276 131356 78328
rect 122288 78208 122340 78260
rect 135444 78208 135496 78260
rect 121276 78140 121328 78192
rect 133696 78140 133748 78192
rect 106924 78072 106976 78124
rect 125232 78072 125284 78124
rect 132316 78072 132368 78124
rect 149980 78276 150032 78328
rect 152464 78276 152516 78328
rect 162308 78276 162360 78328
rect 163136 78276 163188 78328
rect 165528 78276 165580 78328
rect 168564 78276 168616 78328
rect 169392 78276 169444 78328
rect 169668 78276 169720 78328
rect 188712 78276 188764 78328
rect 138940 78208 138992 78260
rect 142252 78208 142304 78260
rect 148876 78208 148928 78260
rect 158168 78208 158220 78260
rect 161204 78208 161256 78260
rect 157248 78140 157300 78192
rect 165988 78140 166040 78192
rect 167276 78208 167328 78260
rect 177396 78208 177448 78260
rect 181812 78208 181864 78260
rect 169484 78140 169536 78192
rect 172980 78140 173032 78192
rect 174728 78140 174780 78192
rect 174820 78140 174872 78192
rect 175004 78140 175056 78192
rect 189724 78140 189776 78192
rect 195244 78140 195296 78192
rect 107476 78004 107528 78056
rect 128452 78004 128504 78056
rect 129004 78004 129056 78056
rect 134248 78004 134300 78056
rect 136732 78004 136784 78056
rect 148784 78072 148836 78124
rect 153384 78072 153436 78124
rect 154120 78072 154172 78124
rect 158168 78072 158220 78124
rect 158812 78072 158864 78124
rect 160376 78072 160428 78124
rect 166172 78072 166224 78124
rect 167460 78072 167512 78124
rect 182088 78072 182140 78124
rect 182916 78072 182968 78124
rect 196808 78072 196860 78124
rect 103980 77936 104032 77988
rect 135904 77936 135956 77988
rect 155684 78004 155736 78056
rect 157892 78004 157944 78056
rect 169668 78004 169720 78056
rect 170496 78004 170548 78056
rect 180524 78004 180576 78056
rect 180708 78004 180760 78056
rect 204996 78004 205048 78056
rect 148324 77936 148376 77988
rect 148968 77936 149020 77988
rect 156512 77936 156564 77988
rect 169300 77936 169352 77988
rect 180340 77936 180392 77988
rect 206376 77936 206428 77988
rect 137376 77868 137428 77920
rect 140504 77868 140556 77920
rect 137928 77800 137980 77852
rect 138388 77800 138440 77852
rect 138572 77800 138624 77852
rect 141424 77800 141476 77852
rect 144368 77800 144420 77852
rect 96252 77732 96304 77784
rect 138848 77732 138900 77784
rect 122012 77664 122064 77716
rect 135076 77664 135128 77716
rect 154028 77868 154080 77920
rect 163228 77868 163280 77920
rect 163964 77868 164016 77920
rect 167276 77868 167328 77920
rect 167552 77868 167604 77920
rect 170956 77868 171008 77920
rect 173532 77868 173584 77920
rect 182824 77868 182876 77920
rect 195612 77868 195664 77920
rect 147772 77800 147824 77852
rect 148600 77800 148652 77852
rect 157708 77732 157760 77784
rect 213000 77732 213052 77784
rect 165804 77664 165856 77716
rect 166356 77664 166408 77716
rect 167920 77664 167972 77716
rect 169024 77664 169076 77716
rect 170312 77664 170364 77716
rect 189908 77664 189960 77716
rect 99104 77528 99156 77580
rect 138572 77596 138624 77648
rect 140320 77596 140372 77648
rect 139952 77528 140004 77580
rect 140596 77528 140648 77580
rect 144828 77528 144880 77580
rect 138756 77460 138808 77512
rect 146300 77460 146352 77512
rect 134156 77324 134208 77376
rect 134892 77324 134944 77376
rect 132132 77256 132184 77308
rect 139124 77256 139176 77308
rect 163596 77596 163648 77648
rect 170956 77596 171008 77648
rect 147772 77528 147824 77580
rect 148692 77528 148744 77580
rect 165068 77460 165120 77512
rect 172520 77460 172572 77512
rect 156880 77256 156932 77308
rect 159456 77256 159508 77308
rect 163872 77256 163924 77308
rect 2780 77188 2832 77240
rect 4804 77188 4856 77240
rect 120080 77188 120132 77240
rect 142344 77188 142396 77240
rect 158628 77188 158680 77240
rect 160560 77188 160612 77240
rect 176108 77188 176160 77240
rect 200488 77188 200540 77240
rect 115296 77120 115348 77172
rect 140044 77120 140096 77172
rect 140228 77120 140280 77172
rect 152924 77120 152976 77172
rect 215576 77120 215628 77172
rect 140412 77052 140464 77104
rect 141700 77052 141752 77104
rect 143080 77052 143132 77104
rect 159272 77052 159324 77104
rect 159456 77052 159508 77104
rect 172428 77052 172480 77104
rect 211896 77052 211948 77104
rect 117780 76984 117832 77036
rect 166540 76984 166592 77036
rect 173624 76984 173676 77036
rect 211804 76984 211856 77036
rect 115848 76916 115900 76968
rect 142620 76916 142672 76968
rect 156052 76916 156104 76968
rect 157708 76916 157760 76968
rect 175372 76916 175424 76968
rect 218428 76916 218480 76968
rect 114100 76848 114152 76900
rect 146116 76848 146168 76900
rect 156420 76848 156472 76900
rect 158720 76848 158772 76900
rect 192484 76848 192536 76900
rect 113732 76780 113784 76832
rect 147588 76780 147640 76832
rect 172796 76780 172848 76832
rect 208952 76780 209004 76832
rect 118332 76712 118384 76764
rect 149244 76712 149296 76764
rect 119344 76644 119396 76696
rect 149612 76644 149664 76696
rect 94964 76576 95016 76628
rect 129648 76576 129700 76628
rect 135628 76576 135680 76628
rect 136088 76576 136140 76628
rect 139584 76576 139636 76628
rect 139860 76576 139912 76628
rect 141332 76576 141384 76628
rect 141700 76576 141752 76628
rect 142620 76576 142672 76628
rect 145012 76576 145064 76628
rect 153752 76576 153804 76628
rect 154488 76576 154540 76628
rect 154672 76576 154724 76628
rect 154856 76576 154908 76628
rect 156512 76576 156564 76628
rect 156972 76576 157024 76628
rect 67640 76508 67692 76560
rect 115204 76508 115256 76560
rect 115848 76508 115900 76560
rect 135536 76508 135588 76560
rect 136364 76508 136416 76560
rect 177488 76712 177540 76764
rect 209964 76712 210016 76764
rect 168472 76644 168524 76696
rect 203340 76644 203392 76696
rect 165712 76576 165764 76628
rect 176476 76576 176528 76628
rect 179788 76576 179840 76628
rect 203064 76576 203116 76628
rect 289820 76508 289872 76560
rect 102140 76440 102192 76492
rect 133144 76440 133196 76492
rect 141056 76440 141108 76492
rect 141792 76440 141844 76492
rect 155316 76440 155368 76492
rect 158536 76440 158588 76492
rect 165712 76440 165764 76492
rect 166816 76440 166868 76492
rect 119160 76372 119212 76424
rect 156420 76372 156472 76424
rect 165528 76372 165580 76424
rect 204812 76372 204864 76424
rect 94688 76304 94740 76356
rect 163504 76304 163556 76356
rect 113640 76236 113692 76288
rect 166448 76236 166500 76288
rect 180340 76304 180392 76356
rect 170036 76236 170088 76288
rect 180708 76236 180760 76288
rect 135720 76168 135772 76220
rect 136456 76168 136508 76220
rect 140964 76168 141016 76220
rect 141608 76168 141660 76220
rect 155132 76168 155184 76220
rect 155592 76168 155644 76220
rect 156420 76168 156472 76220
rect 156604 76168 156656 76220
rect 158260 76168 158312 76220
rect 158720 76168 158772 76220
rect 159088 76168 159140 76220
rect 159364 76168 159416 76220
rect 166264 76168 166316 76220
rect 166908 76168 166960 76220
rect 132684 76100 132736 76152
rect 132868 76100 132920 76152
rect 136180 76100 136232 76152
rect 136548 76100 136600 76152
rect 154948 76100 155000 76152
rect 155408 76100 155460 76152
rect 156236 76100 156288 76152
rect 157340 76100 157392 76152
rect 175188 76100 175240 76152
rect 177948 76100 178000 76152
rect 135352 76032 135404 76084
rect 136456 76032 136508 76084
rect 136824 76032 136876 76084
rect 137284 76032 137336 76084
rect 138020 76032 138072 76084
rect 139032 76032 139084 76084
rect 158996 76032 159048 76084
rect 159364 76032 159416 76084
rect 161756 76032 161808 76084
rect 166264 76032 166316 76084
rect 171232 76032 171284 76084
rect 171876 76032 171928 76084
rect 132868 75964 132920 76016
rect 133880 75964 133932 76016
rect 134064 75964 134116 76016
rect 134432 75964 134484 76016
rect 138480 75964 138532 76016
rect 139124 75964 139176 76016
rect 151084 75964 151136 76016
rect 151360 75964 151412 76016
rect 170680 75964 170732 76016
rect 172060 75964 172112 76016
rect 130384 75896 130436 75948
rect 154304 75896 154356 75948
rect 158996 75896 159048 75948
rect 159272 75896 159324 75948
rect 159916 75896 159968 75948
rect 160560 75896 160612 75948
rect 161756 75896 161808 75948
rect 162124 75896 162176 75948
rect 168472 75896 168524 75948
rect 168840 75896 168892 75948
rect 169944 75896 169996 75948
rect 170128 75896 170180 75948
rect 171324 75896 171376 75948
rect 171692 75896 171744 75948
rect 173348 75896 173400 75948
rect 173716 75896 173768 75948
rect 176752 75896 176804 75948
rect 177672 75896 177724 75948
rect 100392 75828 100444 75880
rect 102140 75828 102192 75880
rect 97356 75760 97408 75812
rect 150164 75828 150216 75880
rect 151084 75828 151136 75880
rect 151636 75828 151688 75880
rect 160284 75828 160336 75880
rect 160836 75828 160888 75880
rect 168748 75828 168800 75880
rect 171784 75828 171836 75880
rect 172244 75828 172296 75880
rect 191932 75828 191984 75880
rect 129648 75760 129700 75812
rect 152832 75760 152884 75812
rect 169852 75760 169904 75812
rect 170864 75760 170916 75812
rect 171600 75760 171652 75812
rect 192944 75760 192996 75812
rect 117320 75692 117372 75744
rect 121092 75692 121144 75744
rect 155776 75692 155828 75744
rect 175556 75692 175608 75744
rect 215392 75692 215444 75744
rect 215852 75692 215904 75744
rect 117044 75624 117096 75676
rect 149244 75624 149296 75676
rect 150164 75624 150216 75676
rect 175832 75624 175884 75676
rect 215484 75624 215536 75676
rect 112812 75556 112864 75608
rect 145932 75556 145984 75608
rect 170772 75556 170824 75608
rect 208492 75556 208544 75608
rect 103244 75488 103296 75540
rect 36544 75216 36596 75268
rect 135260 75488 135312 75540
rect 114376 75420 114428 75472
rect 139952 75420 140004 75472
rect 116952 75352 117004 75404
rect 146668 75488 146720 75540
rect 158260 75488 158312 75540
rect 160652 75488 160704 75540
rect 195152 75488 195204 75540
rect 142252 75420 142304 75472
rect 146208 75420 146260 75472
rect 156052 75420 156104 75472
rect 157064 75420 157116 75472
rect 174544 75420 174596 75472
rect 208584 75420 208636 75472
rect 117872 75284 117924 75336
rect 145104 75352 145156 75404
rect 146392 75352 146444 75404
rect 146852 75352 146904 75404
rect 140872 75284 140924 75336
rect 141976 75284 142028 75336
rect 142344 75284 142396 75336
rect 142896 75284 142948 75336
rect 142988 75284 143040 75336
rect 134248 75216 134300 75268
rect 134800 75216 134852 75268
rect 137008 75216 137060 75268
rect 137652 75216 137704 75268
rect 139952 75216 140004 75268
rect 142252 75216 142304 75268
rect 142620 75216 142672 75268
rect 142804 75216 142856 75268
rect 143908 75216 143960 75268
rect 144276 75216 144328 75268
rect 164240 75216 164292 75268
rect 164608 75216 164660 75268
rect 78680 75148 78732 75200
rect 108856 75080 108908 75132
rect 108488 75012 108540 75064
rect 132132 75012 132184 75064
rect 134156 75012 134208 75064
rect 134524 75012 134576 75064
rect 141056 75080 141108 75132
rect 141884 75080 141936 75132
rect 142528 75012 142580 75064
rect 142988 75012 143040 75064
rect 148140 75148 148192 75200
rect 148324 75148 148376 75200
rect 164332 75148 164384 75200
rect 165344 75148 165396 75200
rect 163412 75080 163464 75132
rect 169208 75352 169260 75404
rect 201776 75352 201828 75404
rect 202788 75352 202840 75404
rect 180524 75284 180576 75336
rect 210240 75284 210292 75336
rect 167184 75216 167236 75268
rect 167736 75216 167788 75268
rect 174084 75216 174136 75268
rect 174360 75216 174412 75268
rect 202788 75216 202840 75268
rect 281540 75216 281592 75268
rect 167092 75148 167144 75200
rect 168288 75148 168340 75200
rect 181444 75148 181496 75200
rect 214104 75148 214156 75200
rect 215392 75148 215444 75200
rect 525800 75148 525852 75200
rect 158260 75012 158312 75064
rect 164240 75012 164292 75064
rect 165160 75012 165212 75064
rect 174544 75080 174596 75132
rect 177948 75080 178000 75132
rect 207296 75080 207348 75132
rect 214656 75012 214708 75064
rect 120356 74944 120408 74996
rect 142436 74944 142488 74996
rect 142804 74944 142856 74996
rect 157156 74944 157208 74996
rect 214748 74944 214800 74996
rect 149704 74876 149756 74928
rect 179972 74876 180024 74928
rect 161296 74808 161348 74860
rect 181812 74808 181864 74860
rect 167184 74740 167236 74792
rect 168104 74740 168156 74792
rect 153936 74604 153988 74656
rect 154212 74604 154264 74656
rect 107292 74468 107344 74520
rect 132408 74468 132460 74520
rect 169300 74468 169352 74520
rect 191012 74468 191064 74520
rect 127532 74400 127584 74452
rect 147772 74400 147824 74452
rect 175740 74400 175792 74452
rect 211712 74400 211764 74452
rect 120540 74332 120592 74384
rect 158628 74332 158680 74384
rect 162308 74332 162360 74384
rect 196532 74332 196584 74384
rect 109776 74264 109828 74316
rect 143540 74264 143592 74316
rect 159456 74264 159508 74316
rect 192300 74264 192352 74316
rect 114744 74196 114796 74248
rect 147680 74196 147732 74248
rect 166632 74196 166684 74248
rect 197452 74196 197504 74248
rect 119988 74128 120040 74180
rect 152372 74128 152424 74180
rect 165620 74128 165672 74180
rect 196164 74128 196216 74180
rect 113916 74060 113968 74112
rect 145748 74060 145800 74112
rect 163872 74060 163924 74112
rect 193864 74060 193916 74112
rect 119528 73992 119580 74044
rect 151452 73992 151504 74044
rect 159732 73992 159784 74044
rect 193588 73992 193640 74044
rect 115388 73924 115440 73976
rect 145288 73924 145340 73976
rect 172520 73924 172572 73976
rect 199292 73924 199344 73976
rect 114008 73856 114060 73908
rect 142160 73856 142212 73908
rect 162676 73856 162728 73908
rect 182180 73856 182232 73908
rect 13084 73788 13136 73840
rect 119528 73788 119580 73840
rect 143540 73788 143592 73840
rect 144184 73788 144236 73840
rect 274640 73788 274692 73840
rect 107476 73720 107528 73772
rect 132040 73720 132092 73772
rect 164700 73720 164752 73772
rect 202972 73720 203024 73772
rect 94780 73652 94832 73704
rect 148876 73652 148928 73704
rect 165988 73652 166040 73704
rect 190736 73652 190788 73704
rect 109592 73584 109644 73636
rect 148048 73584 148100 73636
rect 182088 73584 182140 73636
rect 201684 73584 201736 73636
rect 105544 73516 105596 73568
rect 131212 73516 131264 73568
rect 3148 73108 3200 73160
rect 111800 73108 111852 73160
rect 123576 73108 123628 73160
rect 129280 73108 129332 73160
rect 152096 73108 152148 73160
rect 158168 73108 158220 73160
rect 158628 73108 158680 73160
rect 182180 73108 182232 73160
rect 183468 73108 183520 73160
rect 193680 73108 193732 73160
rect 131212 73040 131264 73092
rect 132316 73040 132368 73092
rect 138940 73040 138992 73092
rect 143632 73040 143684 73092
rect 144092 73040 144144 73092
rect 144460 73040 144512 73092
rect 172336 73040 172388 73092
rect 203800 73040 203852 73092
rect 112720 72972 112772 73024
rect 138756 72972 138808 73024
rect 142988 72972 143040 73024
rect 143172 72972 143224 73024
rect 166264 72972 166316 73024
rect 196716 72972 196768 73024
rect 126336 72904 126388 72956
rect 150808 72904 150860 72956
rect 156788 72904 156840 72956
rect 190920 72904 190972 72956
rect 191748 72904 191800 72956
rect 101956 72836 102008 72888
rect 106280 72836 106332 72888
rect 107476 72836 107528 72888
rect 118516 72836 118568 72888
rect 151912 72836 151964 72888
rect 162584 72836 162636 72888
rect 194692 72836 194744 72888
rect 119068 72768 119120 72820
rect 153292 72768 153344 72820
rect 162768 72768 162820 72820
rect 195980 72768 196032 72820
rect 113456 72700 113508 72752
rect 147864 72700 147916 72752
rect 156512 72700 156564 72752
rect 156788 72700 156840 72752
rect 190460 72700 190512 72752
rect 111524 72632 111576 72684
rect 144460 72632 144512 72684
rect 158352 72632 158404 72684
rect 189356 72632 189408 72684
rect 110236 72564 110288 72616
rect 142988 72564 143040 72616
rect 175648 72564 175700 72616
rect 204444 72564 204496 72616
rect 119712 72496 119764 72548
rect 151820 72496 151872 72548
rect 169484 72496 169536 72548
rect 194600 72496 194652 72548
rect 54484 72428 54536 72480
rect 100300 72428 100352 72480
rect 134984 72428 135036 72480
rect 145196 72428 145248 72480
rect 185584 72428 185636 72480
rect 191748 72428 191800 72480
rect 255320 72428 255372 72480
rect 98644 72360 98696 72412
rect 133788 72360 133840 72412
rect 158628 72360 158680 72412
rect 192392 72360 192444 72412
rect 111800 72292 111852 72344
rect 112628 72292 112680 72344
rect 147496 72292 147548 72344
rect 153844 72292 153896 72344
rect 218060 72292 218112 72344
rect 94596 72224 94648 72276
rect 157616 72224 157668 72276
rect 153936 72020 153988 72072
rect 154212 72020 154264 72072
rect 108580 71680 108632 71732
rect 143356 71680 143408 71732
rect 143724 71680 143776 71732
rect 144184 71680 144236 71732
rect 173808 71680 173860 71732
rect 174912 71680 174964 71732
rect 175280 71680 175332 71732
rect 176108 71680 176160 71732
rect 114836 71612 114888 71664
rect 149152 71612 149204 71664
rect 149888 71612 149940 71664
rect 169392 71612 169444 71664
rect 210148 71680 210200 71732
rect 176568 71612 176620 71664
rect 215300 71612 215352 71664
rect 119896 71544 119948 71596
rect 153844 71544 153896 71596
rect 171416 71544 171468 71596
rect 206008 71544 206060 71596
rect 207112 71544 207164 71596
rect 207296 71544 207348 71596
rect 126244 71476 126296 71528
rect 151084 71476 151136 71528
rect 170496 71476 170548 71528
rect 204260 71476 204312 71528
rect 116676 71408 116728 71460
rect 149796 71408 149848 71460
rect 165436 71408 165488 71460
rect 197912 71408 197964 71460
rect 110788 71340 110840 71392
rect 143724 71340 143776 71392
rect 174728 71340 174780 71392
rect 207112 71340 207164 71392
rect 110972 71272 111024 71324
rect 143540 71272 143592 71324
rect 147036 71272 147088 71324
rect 171784 71272 171836 71324
rect 203156 71272 203208 71324
rect 110696 71204 110748 71256
rect 144368 71204 144420 71256
rect 173440 71204 173492 71256
rect 201684 71204 201736 71256
rect 202144 71204 202196 71256
rect 117688 71136 117740 71188
rect 149520 71136 149572 71188
rect 171508 71136 171560 71188
rect 199752 71136 199804 71188
rect 133696 71068 133748 71120
rect 265624 71068 265676 71120
rect 4804 71000 4856 71052
rect 156788 71000 156840 71052
rect 164792 71000 164844 71052
rect 165344 71000 165396 71052
rect 176108 71000 176160 71052
rect 199568 71000 199620 71052
rect 215300 71000 215352 71052
rect 484400 71000 484452 71052
rect 111432 70932 111484 70984
rect 140596 70932 140648 70984
rect 177028 70932 177080 70984
rect 196348 70932 196400 70984
rect 101772 70864 101824 70916
rect 136548 70864 136600 70916
rect 156420 70864 156472 70916
rect 187056 70864 187108 70916
rect 125600 70388 125652 70440
rect 173808 70388 173860 70440
rect 111616 70320 111668 70372
rect 145380 70320 145432 70372
rect 145564 70320 145616 70372
rect 172612 70320 172664 70372
rect 193404 70320 193456 70372
rect 120724 70252 120776 70304
rect 154672 70252 154724 70304
rect 165896 70252 165948 70304
rect 207756 70252 207808 70304
rect 114284 70184 114336 70236
rect 146852 70184 146904 70236
rect 176752 70184 176804 70236
rect 212908 70184 212960 70236
rect 116768 70116 116820 70168
rect 151360 70116 151412 70168
rect 166080 70116 166132 70168
rect 200212 70116 200264 70168
rect 120632 70048 120684 70100
rect 152004 70048 152056 70100
rect 172060 70048 172112 70100
rect 205640 70048 205692 70100
rect 118240 69980 118292 70032
rect 150716 69980 150768 70032
rect 174176 69980 174228 70032
rect 207388 69980 207440 70032
rect 207664 69980 207716 70032
rect 115572 69912 115624 69964
rect 148600 69912 148652 69964
rect 167828 69912 167880 69964
rect 201500 69912 201552 69964
rect 112904 69844 112956 69896
rect 145472 69844 145524 69896
rect 171968 69844 172020 69896
rect 204260 69844 204312 69896
rect 115848 69776 115900 69828
rect 148232 69776 148284 69828
rect 173348 69776 173400 69828
rect 205640 69776 205692 69828
rect 64144 69708 64196 69760
rect 98736 69708 98788 69760
rect 132960 69708 133012 69760
rect 142804 69708 142856 69760
rect 300860 69708 300912 69760
rect 43444 69640 43496 69692
rect 115664 69640 115716 69692
rect 115848 69640 115900 69692
rect 143448 69640 143500 69692
rect 173900 69640 173952 69692
rect 176844 69640 176896 69692
rect 207296 69640 207348 69692
rect 207388 69640 207440 69692
rect 407120 69640 407172 69692
rect 109684 69572 109736 69624
rect 137376 69572 137428 69624
rect 167644 69572 167696 69624
rect 197820 69572 197872 69624
rect 99288 69504 99340 69556
rect 132776 69504 132828 69556
rect 156604 69504 156656 69556
rect 218336 69504 218388 69556
rect 166080 69028 166132 69080
rect 166264 69028 166316 69080
rect 97908 68960 97960 69012
rect 131120 68960 131172 69012
rect 152740 68960 152792 69012
rect 216128 68960 216180 69012
rect 579988 68960 580040 69012
rect 3148 68892 3200 68944
rect 111892 68892 111944 68944
rect 121736 68892 121788 68944
rect 141240 68892 141292 68944
rect 160468 68892 160520 68944
rect 182824 68892 182876 68944
rect 95056 68824 95108 68876
rect 155316 68824 155368 68876
rect 171876 68824 171928 68876
rect 196440 68824 196492 68876
rect 122196 68756 122248 68808
rect 122840 68756 122892 68808
rect 146576 68756 146628 68808
rect 161388 68756 161440 68808
rect 194876 68756 194928 68808
rect 104808 68688 104860 68740
rect 138664 68688 138716 68740
rect 157524 68688 157576 68740
rect 191840 68688 191892 68740
rect 105912 68620 105964 68672
rect 139492 68620 139544 68672
rect 161940 68620 161992 68672
rect 162768 68620 162820 68672
rect 101864 68552 101916 68604
rect 136364 68552 136416 68604
rect 107016 68484 107068 68536
rect 139860 68484 139912 68536
rect 160008 68484 160060 68536
rect 193496 68620 193548 68672
rect 110144 68416 110196 68468
rect 141424 68416 141476 68468
rect 161296 68416 161348 68468
rect 195520 68552 195572 68604
rect 171968 68484 172020 68536
rect 196900 68484 196952 68536
rect 107200 68348 107252 68400
rect 135628 68348 135680 68400
rect 159180 68348 159232 68400
rect 193772 68416 193824 68468
rect 172060 68348 172112 68400
rect 199660 68348 199712 68400
rect 134616 68280 134668 68332
rect 211804 68280 211856 68332
rect 111708 68212 111760 68264
rect 152556 68212 152608 68264
rect 168932 68212 168984 68264
rect 190460 68212 190512 68264
rect 203616 68212 203668 68264
rect 111892 68144 111944 68196
rect 113088 68144 113140 68196
rect 146484 68144 146536 68196
rect 162308 68144 162360 68196
rect 182916 68144 182968 68196
rect 103060 68076 103112 68128
rect 138388 68076 138440 68128
rect 160376 68076 160428 68128
rect 161388 68076 161440 68128
rect 168104 68076 168156 68128
rect 202052 68076 202104 68128
rect 107568 68008 107620 68060
rect 135536 68008 135588 68060
rect 158444 68008 158496 68060
rect 160468 68008 160520 68060
rect 162768 68008 162820 68060
rect 171968 68008 172020 68060
rect 161848 67940 161900 67992
rect 171876 67940 171928 67992
rect 160560 67872 160612 67924
rect 161296 67872 161348 67924
rect 159088 67600 159140 67652
rect 160008 67600 160060 67652
rect 167368 67600 167420 67652
rect 168104 67600 168156 67652
rect 96436 67532 96488 67584
rect 141056 67532 141108 67584
rect 168196 67532 168248 67584
rect 217508 67532 217560 67584
rect 580632 67532 580684 67584
rect 109960 67464 110012 67516
rect 144000 67464 144052 67516
rect 176660 67464 176712 67516
rect 211620 67464 211672 67516
rect 212448 67464 212500 67516
rect 110052 67396 110104 67448
rect 144276 67396 144328 67448
rect 163228 67396 163280 67448
rect 198096 67396 198148 67448
rect 104624 67328 104676 67380
rect 104716 67260 104768 67312
rect 135260 67260 135312 67312
rect 135444 67328 135496 67380
rect 136088 67328 136140 67380
rect 137008 67328 137060 67380
rect 137284 67328 137336 67380
rect 138664 67328 138716 67380
rect 139308 67328 139360 67380
rect 139400 67328 139452 67380
rect 140504 67328 140556 67380
rect 174084 67328 174136 67380
rect 208676 67328 208728 67380
rect 138020 67260 138072 67312
rect 160284 67260 160336 67312
rect 194784 67260 194836 67312
rect 108948 67192 109000 67244
rect 142344 67192 142396 67244
rect 142804 67192 142856 67244
rect 164516 67192 164568 67244
rect 199016 67192 199068 67244
rect 110420 67124 110472 67176
rect 112536 67124 112588 67176
rect 147128 67124 147180 67176
rect 164608 67124 164660 67176
rect 199108 67124 199160 67176
rect 26240 66852 26292 66904
rect 103152 66852 103204 66904
rect 137192 67056 137244 67108
rect 138020 67056 138072 67108
rect 138756 67056 138808 67108
rect 163688 67056 163740 67108
rect 164148 67056 164200 67108
rect 197728 67056 197780 67108
rect 104348 66988 104400 67040
rect 137284 66988 137336 67040
rect 170404 66988 170456 67040
rect 204536 66988 204588 67040
rect 107384 66920 107436 66972
rect 135168 66920 135220 66972
rect 135260 66920 135312 66972
rect 138664 66920 138716 66972
rect 166908 66920 166960 66972
rect 200212 66920 200264 66972
rect 212448 66920 212500 66972
rect 236000 66920 236052 66972
rect 116492 66852 116544 66904
rect 148140 66852 148192 66904
rect 148324 66852 148376 66904
rect 150164 66852 150216 66904
rect 503720 66852 503772 66904
rect 103428 66784 103480 66836
rect 134340 66784 134392 66836
rect 108764 66716 108816 66768
rect 139400 66716 139452 66768
rect 106096 66648 106148 66700
rect 135444 66648 135496 66700
rect 135168 66580 135220 66632
rect 140688 66580 140740 66632
rect 170404 66308 170456 66360
rect 170956 66308 171008 66360
rect 120816 66172 120868 66224
rect 141148 66172 141200 66224
rect 346400 66240 346452 66292
rect 142620 66172 142672 66224
rect 142896 66172 142948 66224
rect 158904 66172 158956 66224
rect 219808 66172 219860 66224
rect 102784 66104 102836 66156
rect 142712 66104 142764 66156
rect 143448 66104 143500 66156
rect 156328 66104 156380 66156
rect 216680 66104 216732 66156
rect 116216 66036 116268 66088
rect 155592 66036 155644 66088
rect 170036 66036 170088 66088
rect 209780 66036 209832 66088
rect 117228 65968 117280 66020
rect 153384 65968 153436 66020
rect 164424 65968 164476 66020
rect 203248 65968 203300 66020
rect 100024 65900 100076 65952
rect 134892 65900 134944 65952
rect 158076 65900 158128 65952
rect 192116 65900 192168 65952
rect 193128 65900 193180 65952
rect 101312 65832 101364 65884
rect 136456 65832 136508 65884
rect 146944 65832 146996 65884
rect 173808 65832 173860 65884
rect 208400 65832 208452 65884
rect 99932 65764 99984 65816
rect 133052 65764 133104 65816
rect 153936 65764 153988 65816
rect 188344 65764 188396 65816
rect 105360 65696 105412 65748
rect 138204 65696 138256 65748
rect 167184 65696 167236 65748
rect 168288 65696 168340 65748
rect 200672 65696 200724 65748
rect 102048 65628 102100 65680
rect 134156 65628 134208 65680
rect 134892 65628 134944 65680
rect 135904 65628 135956 65680
rect 161756 65628 161808 65680
rect 189448 65628 189500 65680
rect 193128 65628 193180 65680
rect 216680 65628 216732 65680
rect 35164 65492 35216 65544
rect 118424 65492 118476 65544
rect 151268 65560 151320 65612
rect 167276 65560 167328 65612
rect 171140 65560 171192 65612
rect 201960 65560 202012 65612
rect 128452 65492 128504 65544
rect 129004 65492 129056 65544
rect 143448 65492 143500 65544
rect 438860 65492 438912 65544
rect 99840 65424 99892 65476
rect 139584 65424 139636 65476
rect 112168 65356 112220 65408
rect 132500 65356 132552 65408
rect 134156 65356 134208 65408
rect 134708 65356 134760 65408
rect 95148 65288 95200 65340
rect 160192 65288 160244 65340
rect 121828 65220 121880 65272
rect 142896 65220 142948 65272
rect 3148 64812 3200 64864
rect 158444 64812 158496 64864
rect 169852 64812 169904 64864
rect 171048 64812 171100 64864
rect 171232 64812 171284 64864
rect 171876 64812 171928 64864
rect 175464 64812 175516 64864
rect 175924 64812 175976 64864
rect 212540 64812 212592 64864
rect 96344 64744 96396 64796
rect 146668 64744 146720 64796
rect 169944 64744 169996 64796
rect 205732 64744 205784 64796
rect 118608 64676 118660 64728
rect 153752 64676 153804 64728
rect 165804 64676 165856 64728
rect 200856 64676 200908 64728
rect 100576 64608 100628 64660
rect 134616 64608 134668 64660
rect 173992 64608 174044 64660
rect 175188 64608 175240 64660
rect 208768 64608 208820 64660
rect 106188 64540 106240 64592
rect 140044 64540 140096 64592
rect 171876 64540 171928 64592
rect 205916 64540 205968 64592
rect 100668 64472 100720 64524
rect 132868 64472 132920 64524
rect 133788 64472 133840 64524
rect 173256 64472 173308 64524
rect 173808 64472 173860 64524
rect 207020 64472 207072 64524
rect 104256 64404 104308 64456
rect 136824 64404 136876 64456
rect 161664 64404 161716 64456
rect 196072 64404 196124 64456
rect 122104 64336 122156 64388
rect 154120 64336 154172 64388
rect 171048 64336 171100 64388
rect 203892 64336 203944 64388
rect 128360 64268 128412 64320
rect 207572 64268 207624 64320
rect 106004 64200 106056 64252
rect 137836 64200 137888 64252
rect 144000 64200 144052 64252
rect 278780 64200 278832 64252
rect 136824 64132 136876 64184
rect 144920 64132 144972 64184
rect 154856 64132 154908 64184
rect 189080 64132 189132 64184
rect 488540 64132 488592 64184
rect 162860 64064 162912 64116
rect 163044 64064 163096 64116
rect 191288 64064 191340 64116
rect 165436 63996 165488 64048
rect 189264 63996 189316 64048
rect 157708 63928 157760 63980
rect 189080 63928 189132 63980
rect 96160 63452 96212 63504
rect 143080 63452 143132 63504
rect 154028 63452 154080 63504
rect 580356 63452 580408 63504
rect 97172 63384 97224 63436
rect 139124 63384 139176 63436
rect 156880 63384 156932 63436
rect 580540 63384 580592 63436
rect 100484 63316 100536 63368
rect 141424 63316 141476 63368
rect 156236 63316 156288 63368
rect 215668 63316 215720 63368
rect 96528 63248 96580 63300
rect 134248 63248 134300 63300
rect 161480 63248 161532 63300
rect 219532 63248 219584 63300
rect 162492 63180 162544 63232
rect 210056 63180 210108 63232
rect 167920 63112 167972 63164
rect 210516 63112 210568 63164
rect 164332 63044 164384 63096
rect 165528 63044 165580 63096
rect 206284 63044 206336 63096
rect 167092 62976 167144 63028
rect 208860 62976 208912 63028
rect 165712 62908 165764 62960
rect 166908 62908 166960 62960
rect 207204 62908 207256 62960
rect 31024 62840 31076 62892
rect 162860 62840 162912 62892
rect 168564 62840 168616 62892
rect 182180 62840 182232 62892
rect 219440 62840 219492 62892
rect 142988 62772 143040 62824
rect 430580 62772 430632 62824
rect 167736 62704 167788 62756
rect 202236 62704 202288 62756
rect 134248 62092 134300 62144
rect 134800 62092 134852 62144
rect 138848 62092 138900 62144
rect 139124 62092 139176 62144
rect 158720 62024 158772 62076
rect 193220 62024 193272 62076
rect 194508 62024 194560 62076
rect 155868 61956 155920 62008
rect 186320 61956 186372 62008
rect 161204 61888 161256 61940
rect 190552 61888 190604 61940
rect 137836 61412 137888 61464
rect 385040 61412 385092 61464
rect 22744 61344 22796 61396
rect 174820 61344 174872 61396
rect 194508 61344 194560 61396
rect 558184 61344 558236 61396
rect 160100 61208 160152 61260
rect 161204 61208 161256 61260
rect 96068 60664 96120 60716
rect 139952 60664 140004 60716
rect 168472 60664 168524 60716
rect 219716 60664 219768 60716
rect 220728 60664 220780 60716
rect 93124 60052 93176 60104
rect 167092 60052 167144 60104
rect 220728 60052 220780 60104
rect 404360 60052 404412 60104
rect 48320 59984 48372 60036
rect 96068 59984 96120 60036
rect 144460 59984 144512 60036
rect 342260 59984 342312 60036
rect 169668 59304 169720 59356
rect 203524 59304 203576 59356
rect 204168 59304 204220 59356
rect 166172 59236 166224 59288
rect 201132 59236 201184 59288
rect 201408 59236 201460 59288
rect 201408 58692 201460 58744
rect 251180 58692 251232 58744
rect 95240 58624 95292 58676
rect 166264 58624 166316 58676
rect 204168 58624 204220 58676
rect 510620 58624 510672 58676
rect 169760 57876 169812 57928
rect 204904 57876 204956 57928
rect 155500 57808 155552 57860
rect 189080 57808 189132 57860
rect 189540 57808 189592 57860
rect 204904 57264 204956 57316
rect 231860 57264 231912 57316
rect 6920 57196 6972 57248
rect 160100 57196 160152 57248
rect 189080 57196 189132 57248
rect 560300 57196 560352 57248
rect 3424 56516 3476 56568
rect 97264 56516 97316 56568
rect 155408 56516 155460 56568
rect 214564 56516 214616 56568
rect 17960 55904 18012 55956
rect 176108 55904 176160 55956
rect 214564 55904 214616 55956
rect 376760 55904 376812 55956
rect 133788 55836 133840 55888
rect 538220 55836 538272 55888
rect 101404 55156 101456 55208
rect 135720 55156 135772 55208
rect 162952 55156 163004 55208
rect 198280 55156 198332 55208
rect 145656 54544 145708 54596
rect 224960 54544 225012 54596
rect 13820 54476 13872 54528
rect 101404 54476 101456 54528
rect 198280 54476 198332 54528
rect 400220 54476 400272 54528
rect 105452 53728 105504 53780
rect 138572 53728 138624 53780
rect 141424 53116 141476 53168
rect 205640 53116 205692 53168
rect 3516 53048 3568 53100
rect 105452 53048 105504 53100
rect 149888 53048 149940 53100
rect 469220 53048 469272 53100
rect 3424 52368 3476 52420
rect 110328 52368 110380 52420
rect 138940 52368 138992 52420
rect 164240 52368 164292 52420
rect 219624 52368 219676 52420
rect 220728 52368 220780 52420
rect 149796 51756 149848 51808
rect 309140 51756 309192 51808
rect 220728 51688 220780 51740
rect 563704 51688 563756 51740
rect 164056 51008 164108 51060
rect 197452 51008 197504 51060
rect 149704 50396 149756 50448
rect 305000 50396 305052 50448
rect 197452 50328 197504 50380
rect 543004 50328 543056 50380
rect 3240 49648 3292 49700
rect 162124 49648 162176 49700
rect 183468 49648 183520 49700
rect 580172 49648 580224 49700
rect 140136 48968 140188 49020
rect 374000 48968 374052 49020
rect 156144 48220 156196 48272
rect 190644 48220 190696 48272
rect 191748 48220 191800 48272
rect 191748 47608 191800 47660
rect 369860 47608 369912 47660
rect 137284 47540 137336 47592
rect 442264 47540 442316 47592
rect 156052 46860 156104 46912
rect 215668 46860 215720 46912
rect 216036 46860 216088 46912
rect 215668 46248 215720 46300
rect 396080 46248 396132 46300
rect 134800 46180 134852 46232
rect 324320 46180 324372 46232
rect 3516 45500 3568 45552
rect 22744 45500 22796 45552
rect 147036 45500 147088 45552
rect 579988 45500 580040 45552
rect 144368 43460 144420 43512
rect 354680 43460 354732 43512
rect 140044 43392 140096 43444
rect 456800 43392 456852 43444
rect 134708 42100 134760 42152
rect 242900 42100 242952 42152
rect 161296 42032 161348 42084
rect 521660 42032 521712 42084
rect 3516 41352 3568 41404
rect 122196 41352 122248 41404
rect 185584 41352 185636 41404
rect 580172 41352 580224 41404
rect 148324 40672 148376 40724
rect 193220 40672 193272 40724
rect 161388 39312 161440 39364
rect 578884 39312 578936 39364
rect 164148 37952 164200 38004
rect 331220 37952 331272 38004
rect 137100 37884 137152 37936
rect 389180 37884 389232 37936
rect 3148 37204 3200 37256
rect 128452 37204 128504 37256
rect 155960 37204 156012 37256
rect 197360 37204 197412 37256
rect 580172 37204 580224 37256
rect 165344 35232 165396 35284
rect 247040 35232 247092 35284
rect 153936 35164 153988 35216
rect 499580 35164 499632 35216
rect 168196 33736 168248 33788
rect 423680 33736 423732 33788
rect 158536 33056 158588 33108
rect 580172 33056 580224 33108
rect 3148 32988 3200 33040
rect 177304 32988 177356 33040
rect 168288 31016 168340 31068
rect 495440 31016 495492 31068
rect 162676 29656 162728 29708
rect 357440 29656 357492 29708
rect 133144 29588 133196 29640
rect 507860 29588 507912 29640
rect 3148 28908 3200 28960
rect 147772 28908 147824 28960
rect 170956 28296 171008 28348
rect 296720 28296 296772 28348
rect 144276 28228 144328 28280
rect 571340 28228 571392 28280
rect 175188 26868 175240 26920
rect 480260 26868 480312 26920
rect 167000 26256 167052 26308
rect 171876 26256 171928 26308
rect 173808 25576 173860 25628
rect 262220 25576 262272 25628
rect 155868 25508 155920 25560
rect 575480 25508 575532 25560
rect 3056 24760 3108 24812
rect 35164 24760 35216 24812
rect 184204 24760 184256 24812
rect 580172 24760 580224 24812
rect 171048 22788 171100 22840
rect 350540 22788 350592 22840
rect 138756 22720 138808 22772
rect 392584 22720 392636 22772
rect 144184 21428 144236 21480
rect 320180 21428 320232 21480
rect 138848 21360 138900 21412
rect 434720 21360 434772 21412
rect 3516 20612 3568 20664
rect 139400 20612 139452 20664
rect 180708 20612 180760 20664
rect 580172 20612 580224 20664
rect 160008 18640 160060 18692
rect 361580 18640 361632 18692
rect 134616 18572 134668 18624
rect 454040 18572 454092 18624
rect 153844 17212 153896 17264
rect 465080 17212 465132 17264
rect 3516 16532 3568 16584
rect 131212 16532 131264 16584
rect 165436 16532 165488 16584
rect 580172 16532 580224 16584
rect 151084 14492 151136 14544
rect 316408 14492 316460 14544
rect 166908 14424 166960 14476
rect 549536 14424 549588 14476
rect 142896 13064 142948 13116
rect 477224 13064 477276 13116
rect 3056 12384 3108 12436
rect 130384 12384 130436 12436
rect 182088 12384 182140 12436
rect 580172 12384 580224 12436
rect 137192 10344 137244 10396
rect 176016 10344 176068 10396
rect 142804 10276 142856 10328
rect 418804 10276 418856 10328
rect 160376 9052 160428 9104
rect 175924 9052 175976 9104
rect 145564 8984 145616 9036
rect 340052 8984 340104 9036
rect 134524 8916 134576 8968
rect 530676 8916 530728 8968
rect 2964 8236 3016 8288
rect 13084 8236 13136 8288
rect 152464 8236 152516 8288
rect 580172 8236 580224 8288
rect 165528 7556 165580 7608
rect 461768 7556 461820 7608
rect 162768 6128 162820 6180
rect 473360 6128 473412 6180
rect 543004 5448 543056 5500
rect 580172 5448 580224 5500
rect 152648 4836 152700 4888
rect 171784 4836 171836 4888
rect 38016 4768 38068 4820
rect 116584 4768 116636 4820
rect 158628 4768 158680 4820
rect 542268 4768 542320 4820
rect 148784 4632 148836 4684
rect 151912 4632 151964 4684
rect 3148 4088 3200 4140
rect 54484 4088 54536 4140
rect 34152 3680 34204 3732
rect 36544 3680 36596 3732
rect 174544 3612 174596 3664
rect 186780 3612 186832 3664
rect 20 3544 72 3596
rect 3332 3544 3384 3596
rect 91468 3544 91520 3596
rect 93124 3544 93176 3596
rect 97816 3544 97868 3596
rect 179052 3544 179104 3596
rect 242900 3544 242952 3596
rect 244096 3544 244148 3596
rect 262220 3544 262272 3596
rect 263416 3544 263468 3596
rect 265624 3544 265676 3596
rect 267280 3544 267332 3596
rect 281540 3544 281592 3596
rect 282736 3544 282788 3596
rect 357440 3544 357492 3596
rect 358728 3544 358780 3596
rect 3240 3476 3292 3528
rect 4804 3476 4856 3528
rect 30288 3476 30340 3528
rect 31024 3476 31076 3528
rect 41880 3476 41932 3528
rect 43444 3476 43496 3528
rect 48320 3476 48372 3528
rect 49608 3476 49660 3528
rect 53472 3476 53524 3528
rect 64144 3476 64196 3528
rect 72148 3476 72200 3528
rect 64420 3408 64472 3460
rect 135444 3408 135496 3460
rect 135904 3476 135956 3528
rect 141056 3476 141108 3528
rect 146944 3476 146996 3528
rect 381912 3476 381964 3528
rect 395344 3476 395396 3528
rect 416044 3476 416096 3528
rect 418804 3476 418856 3528
rect 419908 3476 419960 3528
rect 442264 3476 442316 3528
rect 443092 3476 443144 3528
rect 571340 3476 571392 3528
rect 572536 3476 572588 3528
rect 138664 3408 138716 3460
rect 557724 3408 557776 3460
rect 558184 3408 558236 3460
rect 568672 3408 568724 3460
rect 139492 3340 139544 3392
rect 211804 3000 211856 3052
rect 213828 3000 213880 3052
rect 392584 3000 392636 3052
rect 393504 3000 393556 3052
rect 563704 3000 563756 3052
rect 565452 3000 565504 3052
rect 376760 2592 376812 2644
rect 378048 2592 378100 2644
rect 396080 2592 396132 2644
rect 397368 2592 397420 2644
<< metal2 >>
rect 1278 703520 1390 704960
rect 4172 703582 5028 703610
rect 3054 701856 3110 701865
rect 3054 701791 3110 701800
rect 3068 701078 3096 701791
rect 3056 701072 3108 701078
rect 3056 701014 3108 701020
rect 3146 693696 3202 693705
rect 3146 693631 3202 693640
rect 3160 692850 3188 693631
rect 3148 692844 3200 692850
rect 3148 692786 3200 692792
rect 3422 689616 3478 689625
rect 3422 689551 3478 689560
rect 3436 688702 3464 689551
rect 3424 688696 3476 688702
rect 3424 688638 3476 688644
rect 3146 685536 3202 685545
rect 3146 685471 3202 685480
rect 3160 684554 3188 685471
rect 3148 684548 3200 684554
rect 3148 684490 3200 684496
rect 3422 681456 3478 681465
rect 3422 681391 3478 681400
rect 3436 680406 3464 681391
rect 3424 680400 3476 680406
rect 3424 680342 3476 680348
rect 3238 673296 3294 673305
rect 3238 673231 3294 673240
rect 3252 672110 3280 673231
rect 3240 672104 3292 672110
rect 3240 672046 3292 672052
rect 3422 669216 3478 669225
rect 3422 669151 3478 669160
rect 3436 667962 3464 669151
rect 3424 667956 3476 667962
rect 3424 667898 3476 667904
rect 3238 665136 3294 665145
rect 3238 665071 3294 665080
rect 3252 663814 3280 665071
rect 3240 663808 3292 663814
rect 3240 663750 3292 663756
rect 3424 661088 3476 661094
rect 3422 661056 3424 661065
rect 3476 661056 3478 661065
rect 3422 660991 3478 661000
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 645416 3478 645425
rect 3422 645351 3478 645360
rect 3436 644502 3464 645351
rect 3424 644496 3476 644502
rect 3424 644438 3476 644444
rect 3422 629096 3478 629105
rect 3422 629031 3478 629040
rect 3436 627978 3464 629031
rect 3424 627972 3476 627978
rect 3424 627914 3476 627920
rect 3238 625016 3294 625025
rect 3238 624951 3294 624960
rect 3252 623830 3280 624951
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3422 620936 3478 620945
rect 3422 620871 3478 620880
rect 3436 619682 3464 620871
rect 3424 619676 3476 619682
rect 3424 619618 3476 619624
rect 3238 616856 3294 616865
rect 3238 616791 3294 616800
rect 3252 615534 3280 616791
rect 3240 615528 3292 615534
rect 3240 615470 3292 615476
rect 3424 612808 3476 612814
rect 3422 612776 3424 612785
rect 3476 612776 3478 612785
rect 3422 612711 3478 612720
rect 3422 608696 3478 608705
rect 3422 608631 3424 608640
rect 3476 608631 3478 608640
rect 3424 608602 3476 608608
rect 3422 604616 3478 604625
rect 3422 604551 3478 604560
rect 3436 604518 3464 604551
rect 3424 604512 3476 604518
rect 3424 604454 3476 604460
rect 3422 600536 3478 600545
rect 3422 600471 3478 600480
rect 3436 600370 3464 600471
rect 3424 600364 3476 600370
rect 3424 600306 3476 600312
rect 3422 597136 3478 597145
rect 3422 597071 3478 597080
rect 3436 596222 3464 597071
rect 3424 596216 3476 596222
rect 3424 596158 3476 596164
rect 3422 588976 3478 588985
rect 3422 588911 3478 588920
rect 3436 587926 3464 588911
rect 3424 587920 3476 587926
rect 3424 587862 3476 587868
rect 3422 584896 3478 584905
rect 3422 584831 3478 584840
rect 3436 583778 3464 584831
rect 3424 583772 3476 583778
rect 3424 583714 3476 583720
rect 3422 580816 3478 580825
rect 3422 580751 3478 580760
rect 3436 579698 3464 580751
rect 3424 579692 3476 579698
rect 3424 579634 3476 579640
rect 3238 576736 3294 576745
rect 3238 576671 3294 576680
rect 3252 575550 3280 576671
rect 3240 575544 3292 575550
rect 3240 575486 3292 575492
rect 3422 572656 3478 572665
rect 3422 572591 3478 572600
rect 3436 571402 3464 572591
rect 3424 571396 3476 571402
rect 3424 571338 3476 571344
rect 3238 568576 3294 568585
rect 3238 568511 3294 568520
rect 3252 567254 3280 568511
rect 3240 567248 3292 567254
rect 3240 567190 3292 567196
rect 3422 564496 3478 564505
rect 3422 564431 3424 564440
rect 3476 564431 3478 564440
rect 3424 564402 3476 564408
rect 3422 560416 3478 560425
rect 3422 560351 3478 560360
rect 3436 560318 3464 560351
rect 3424 560312 3476 560318
rect 3424 560254 3476 560260
rect 3422 556336 3478 556345
rect 3422 556271 3478 556280
rect 3436 556238 3464 556271
rect 3424 556232 3476 556238
rect 3424 556174 3476 556180
rect 3422 552256 3478 552265
rect 3422 552191 3478 552200
rect 3436 552090 3464 552191
rect 3424 552084 3476 552090
rect 3424 552026 3476 552032
rect 3238 548176 3294 548185
rect 3238 548111 3294 548120
rect 3252 547942 3280 548111
rect 3240 547936 3292 547942
rect 3240 547878 3292 547884
rect 3330 544096 3386 544105
rect 3330 544031 3386 544040
rect 3344 543794 3372 544031
rect 3332 543788 3384 543794
rect 3332 543730 3384 543736
rect 3422 540016 3478 540025
rect 3422 539951 3478 539960
rect 3436 539646 3464 539951
rect 3424 539640 3476 539646
rect 3424 539582 3476 539588
rect 3238 532536 3294 532545
rect 3238 532471 3294 532480
rect 3252 531350 3280 532471
rect 3240 531344 3292 531350
rect 3240 531286 3292 531292
rect 3422 528456 3478 528465
rect 3422 528391 3478 528400
rect 3436 527202 3464 528391
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3238 524376 3294 524385
rect 3238 524311 3294 524320
rect 3252 523054 3280 524311
rect 3240 523048 3292 523054
rect 3240 522990 3292 522996
rect 3424 520328 3476 520334
rect 3422 520296 3424 520305
rect 3476 520296 3478 520305
rect 3422 520231 3478 520240
rect 3422 516216 3478 516225
rect 3422 516151 3424 516160
rect 3476 516151 3478 516160
rect 3424 516122 3476 516128
rect 3422 512136 3478 512145
rect 3422 512071 3478 512080
rect 3436 512038 3464 512071
rect 3424 512032 3476 512038
rect 3424 511974 3476 511980
rect 3422 508056 3478 508065
rect 3422 507991 3478 508000
rect 3436 507890 3464 507991
rect 3424 507884 3476 507890
rect 3424 507826 3476 507832
rect 3238 503976 3294 503985
rect 3238 503911 3294 503920
rect 3252 503742 3280 503911
rect 3240 503736 3292 503742
rect 3240 503678 3292 503684
rect 3330 499896 3386 499905
rect 3330 499831 3386 499840
rect 3344 499594 3372 499831
rect 3332 499588 3384 499594
rect 3332 499530 3384 499536
rect 2870 495816 2926 495825
rect 2870 495751 2926 495760
rect 2884 495514 2912 495751
rect 2872 495508 2924 495514
rect 2872 495450 2924 495456
rect 3422 491736 3478 491745
rect 3422 491671 3478 491680
rect 3436 491366 3464 491671
rect 3424 491360 3476 491366
rect 3424 491302 3476 491308
rect 3422 487656 3478 487665
rect 3422 487591 3478 487600
rect 3436 487218 3464 487591
rect 3424 487212 3476 487218
rect 3424 487154 3476 487160
rect 3514 483576 3570 483585
rect 3514 483511 3570 483520
rect 3528 483070 3556 483511
rect 3516 483064 3568 483070
rect 3516 483006 3568 483012
rect 3422 480176 3478 480185
rect 3422 480111 3478 480120
rect 3436 478922 3464 480111
rect 3424 478916 3476 478922
rect 3424 478858 3476 478864
rect 3238 476096 3294 476105
rect 3238 476031 3294 476040
rect 3252 474774 3280 476031
rect 3240 474768 3292 474774
rect 3240 474710 3292 474716
rect 3424 472048 3476 472054
rect 3422 472016 3424 472025
rect 3476 472016 3478 472025
rect 3422 471951 3478 471960
rect 3422 467936 3478 467945
rect 3422 467871 3424 467880
rect 3476 467871 3478 467880
rect 3424 467842 3476 467848
rect 3422 463856 3478 463865
rect 3422 463791 3478 463800
rect 3436 463758 3464 463791
rect 3424 463752 3476 463758
rect 3424 463694 3476 463700
rect 3422 459776 3478 459785
rect 3422 459711 3478 459720
rect 3436 459610 3464 459711
rect 3424 459604 3476 459610
rect 3424 459546 3476 459552
rect 3238 455696 3294 455705
rect 3238 455631 3294 455640
rect 3252 455462 3280 455631
rect 3240 455456 3292 455462
rect 3240 455398 3292 455404
rect 3330 451616 3386 451625
rect 3330 451551 3386 451560
rect 3344 451314 3372 451551
rect 3332 451308 3384 451314
rect 3332 451250 3384 451256
rect 3422 443456 3478 443465
rect 3422 443391 3478 443400
rect 3436 443018 3464 443391
rect 3424 443012 3476 443018
rect 3424 442954 3476 442960
rect 3422 439376 3478 439385
rect 3422 439311 3478 439320
rect 2870 427136 2926 427145
rect 2870 427071 2926 427080
rect 2884 426494 2912 427071
rect 2872 426488 2924 426494
rect 2872 426430 2924 426436
rect 2962 423056 3018 423065
rect 2962 422991 3018 423000
rect 2976 422346 3004 422991
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 403336 3386 403345
rect 3330 403271 3386 403280
rect 3344 403034 3372 403271
rect 3332 403028 3384 403034
rect 3332 402970 3384 402976
rect 2870 378856 2926 378865
rect 2870 378791 2926 378800
rect 2884 378214 2912 378791
rect 2872 378208 2924 378214
rect 2872 378150 2924 378156
rect 2962 374776 3018 374785
rect 2962 374711 3018 374720
rect 2976 374066 3004 374711
rect 2964 374060 3016 374066
rect 2964 374002 3016 374008
rect 3054 370696 3110 370705
rect 3054 370631 3110 370640
rect 3068 369918 3096 370631
rect 3056 369912 3108 369918
rect 3056 369854 3108 369860
rect 3054 362536 3110 362545
rect 3054 362471 3110 362480
rect 3068 361622 3096 362471
rect 3056 361616 3108 361622
rect 3056 361558 3108 361564
rect 3330 359136 3386 359145
rect 3330 359071 3386 359080
rect 3344 358834 3372 359071
rect 3332 358828 3384 358834
rect 3332 358770 3384 358776
rect 3330 355056 3386 355065
rect 3330 354991 3386 355000
rect 3344 354754 3372 354991
rect 3332 354748 3384 354754
rect 3332 354690 3384 354696
rect 3330 346896 3386 346905
rect 3330 346831 3386 346840
rect 3344 346458 3372 346831
rect 3332 346452 3384 346458
rect 3332 346394 3384 346400
rect 2962 330576 3018 330585
rect 2962 330511 3018 330520
rect 2976 329866 3004 330511
rect 2964 329860 3016 329866
rect 2964 329802 3016 329808
rect 3054 322416 3110 322425
rect 3054 322351 3110 322360
rect 3068 321638 3096 322351
rect 3056 321632 3108 321638
rect 3056 321574 3108 321580
rect 3054 314256 3110 314265
rect 3054 314191 3110 314200
rect 3068 313342 3096 314191
rect 3056 313336 3108 313342
rect 3056 313278 3108 313284
rect 3146 310176 3202 310185
rect 3146 310111 3202 310120
rect 3160 309194 3188 310111
rect 3148 309188 3200 309194
rect 3148 309130 3200 309136
rect 3238 306096 3294 306105
rect 3238 306031 3294 306040
rect 3252 305046 3280 306031
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3146 302016 3202 302025
rect 3146 301951 3202 301960
rect 3160 300898 3188 301951
rect 3148 300892 3200 300898
rect 3148 300834 3200 300840
rect 3330 298616 3386 298625
rect 3330 298551 3386 298560
rect 3344 298178 3372 298551
rect 3332 298172 3384 298178
rect 3332 298114 3384 298120
rect 2870 286376 2926 286385
rect 2870 286311 2926 286320
rect 2884 285734 2912 286311
rect 2872 285728 2924 285734
rect 2872 285670 2924 285676
rect 2962 282296 3018 282305
rect 2962 282231 3018 282240
rect 2976 281586 3004 282231
rect 2964 281580 3016 281586
rect 2964 281522 3016 281528
rect 3054 278216 3110 278225
rect 3054 278151 3110 278160
rect 3068 277438 3096 278151
rect 3056 277432 3108 277438
rect 3056 277374 3108 277380
rect 3054 270056 3110 270065
rect 3054 269991 3110 270000
rect 3068 269142 3096 269991
rect 3056 269136 3108 269142
rect 3056 269078 3108 269084
rect 3146 265976 3202 265985
rect 3146 265911 3202 265920
rect 3160 264994 3188 265911
rect 3148 264988 3200 264994
rect 3148 264930 3200 264936
rect 3054 261896 3110 261905
rect 3054 261831 3110 261840
rect 3068 260982 3096 261831
rect 3056 260976 3108 260982
rect 3056 260918 3108 260924
rect 3238 257816 3294 257825
rect 3238 257751 3294 257760
rect 3252 256766 3280 257751
rect 3240 256760 3292 256766
rect 3240 256702 3292 256708
rect 3146 253736 3202 253745
rect 3146 253671 3202 253680
rect 3160 252618 3188 253671
rect 3148 252612 3200 252618
rect 3148 252554 3200 252560
rect 3330 241496 3386 241505
rect 3330 241431 3386 241440
rect 3344 240174 3372 241431
rect 3332 240168 3384 240174
rect 3332 240110 3384 240116
rect 3330 229936 3386 229945
rect 3330 229871 3386 229880
rect 3344 229158 3372 229871
rect 3332 229152 3384 229158
rect 3332 229094 3384 229100
rect 3054 221776 3110 221785
rect 3054 221711 3110 221720
rect 3068 220862 3096 221711
rect 3056 220856 3108 220862
rect 3056 220798 3108 220804
rect 3146 209536 3202 209545
rect 3146 209471 3202 209480
rect 3160 208418 3188 209471
rect 3148 208412 3200 208418
rect 3148 208354 3200 208360
rect 3146 197296 3202 197305
rect 3146 197231 3202 197240
rect 3160 196654 3188 197231
rect 3148 196648 3200 196654
rect 3148 196590 3200 196596
rect 3436 193866 3464 439311
rect 3514 431216 3570 431225
rect 3514 431151 3570 431160
rect 3528 430642 3556 431151
rect 3516 430636 3568 430642
rect 3516 430578 3568 430584
rect 3514 419656 3570 419665
rect 3514 419591 3570 419600
rect 3528 419558 3556 419591
rect 3516 419552 3568 419558
rect 3516 419494 3568 419500
rect 3514 415576 3570 415585
rect 3514 415511 3570 415520
rect 3528 415478 3556 415511
rect 3516 415472 3568 415478
rect 3516 415414 3568 415420
rect 3514 411496 3570 411505
rect 3514 411431 3570 411440
rect 3528 411330 3556 411431
rect 3516 411324 3568 411330
rect 3516 411266 3568 411272
rect 3514 407416 3570 407425
rect 3514 407351 3570 407360
rect 3528 407182 3556 407351
rect 3516 407176 3568 407182
rect 3516 407118 3568 407124
rect 3514 391096 3570 391105
rect 3514 391031 3570 391040
rect 3528 390590 3556 391031
rect 3516 390584 3568 390590
rect 3516 390526 3568 390532
rect 3514 387016 3570 387025
rect 3514 386951 3570 386960
rect 3528 386442 3556 386951
rect 3516 386436 3568 386442
rect 3516 386378 3568 386384
rect 3514 350976 3570 350985
rect 3514 350911 3570 350920
rect 3528 350606 3556 350911
rect 3516 350600 3568 350606
rect 3516 350542 3568 350548
rect 3514 342816 3570 342825
rect 3514 342751 3570 342760
rect 3528 342310 3556 342751
rect 3516 342304 3568 342310
rect 3516 342246 3568 342252
rect 3514 338736 3570 338745
rect 3514 338671 3570 338680
rect 3528 338162 3556 338671
rect 3516 338156 3568 338162
rect 3516 338098 3568 338104
rect 3514 318336 3570 318345
rect 3514 318271 3570 318280
rect 3528 317490 3556 318271
rect 3516 317484 3568 317490
rect 3516 317426 3568 317432
rect 3514 294536 3570 294545
rect 3514 294471 3570 294480
rect 3528 294030 3556 294471
rect 3516 294024 3568 294030
rect 3516 293966 3568 293972
rect 3514 290456 3570 290465
rect 3514 290391 3570 290400
rect 3528 289882 3556 290391
rect 3516 289876 3568 289882
rect 3516 289818 3568 289824
rect 3514 274136 3570 274145
rect 3514 274071 3570 274080
rect 3528 273290 3556 274071
rect 3516 273284 3568 273290
rect 3516 273226 3568 273232
rect 3514 249656 3570 249665
rect 3514 249591 3570 249600
rect 3528 200802 3556 249591
rect 3606 225856 3662 225865
rect 3606 225791 3662 225800
rect 3620 200870 3648 225791
rect 4066 201376 4122 201385
rect 4066 201311 4122 201320
rect 3608 200864 3660 200870
rect 3608 200806 3660 200812
rect 3516 200796 3568 200802
rect 3516 200738 3568 200744
rect 4080 199442 4108 201311
rect 4068 199436 4120 199442
rect 4068 199378 4120 199384
rect 4172 199345 4200 703582
rect 5000 703474 5028 703582
rect 5142 703520 5254 704960
rect 8312 703582 8892 703610
rect 5184 703474 5212 703520
rect 5000 703446 5212 703474
rect 7564 564460 7616 564466
rect 7564 564402 7616 564408
rect 7576 267034 7604 564402
rect 7564 267028 7616 267034
rect 7564 266970 7616 266976
rect 7564 260908 7616 260914
rect 7564 260850 7616 260856
rect 4158 199336 4214 199345
rect 4158 199271 4214 199280
rect 4804 195288 4856 195294
rect 4804 195230 4856 195236
rect 3424 193860 3476 193866
rect 3424 193802 3476 193808
rect 3422 193216 3478 193225
rect 3422 193151 3478 193160
rect 3436 192506 3464 193151
rect 3424 192500 3476 192506
rect 3424 192442 3476 192448
rect 3422 189136 3478 189145
rect 3422 189071 3424 189080
rect 3476 189071 3478 189080
rect 3424 189042 3476 189048
rect 3424 185156 3476 185162
rect 3424 185098 3476 185104
rect 3436 185065 3464 185098
rect 3422 185056 3478 185065
rect 3422 184991 3478 185000
rect 3422 180976 3478 180985
rect 3422 180911 3478 180920
rect 3436 180878 3464 180911
rect 3424 180872 3476 180878
rect 3424 180814 3476 180820
rect 3330 177576 3386 177585
rect 3330 177511 3386 177520
rect 3344 171134 3372 177511
rect 3422 173496 3478 173505
rect 3422 173431 3478 173440
rect 3436 172582 3464 173431
rect 3424 172576 3476 172582
rect 3424 172518 3476 172524
rect 3344 171106 3464 171134
rect 3146 169416 3202 169425
rect 3146 169351 3202 169360
rect 3160 168434 3188 169351
rect 3148 168428 3200 168434
rect 3148 168370 3200 168376
rect 2780 165368 2832 165374
rect 2778 165336 2780 165345
rect 2832 165336 2834 165345
rect 2778 165271 2834 165280
rect 3436 149138 3464 171106
rect 4816 165374 4844 195230
rect 7576 185162 7604 260850
rect 8312 186114 8340 703582
rect 8864 703474 8892 703582
rect 9006 703520 9118 704960
rect 12452 703582 12756 703610
rect 9048 703474 9076 703520
rect 8864 703446 9076 703474
rect 10324 527196 10376 527202
rect 10324 527138 10376 527144
rect 10336 268462 10364 527138
rect 10324 268456 10376 268462
rect 10324 268398 10376 268404
rect 8944 190528 8996 190534
rect 8944 190470 8996 190476
rect 8300 186108 8352 186114
rect 8300 186050 8352 186056
rect 7564 185156 7616 185162
rect 7564 185098 7616 185104
rect 4804 165368 4856 165374
rect 4804 165310 4856 165316
rect 3516 161424 3568 161430
rect 3516 161366 3568 161372
rect 3528 161265 3556 161366
rect 3514 161256 3570 161265
rect 3514 161191 3570 161200
rect 3514 157176 3570 157185
rect 3514 157111 3570 157120
rect 3528 155990 3556 157111
rect 3516 155984 3568 155990
rect 3516 155926 3568 155932
rect 3514 153096 3570 153105
rect 3514 153031 3570 153040
rect 3528 151842 3556 153031
rect 3516 151836 3568 151842
rect 3516 151778 3568 151784
rect 3436 149110 3556 149138
rect 3424 149048 3476 149054
rect 3422 149016 3424 149025
rect 3476 149016 3478 149025
rect 3422 148951 3478 148960
rect 3424 144968 3476 144974
rect 3422 144936 3424 144945
rect 3476 144936 3478 144945
rect 3528 144906 3556 149110
rect 3422 144871 3478 144880
rect 3516 144900 3568 144906
rect 3516 144842 3568 144848
rect 8956 141370 8984 190470
rect 12452 190233 12480 703582
rect 12728 703474 12756 703582
rect 12870 703520 12982 704960
rect 16090 703520 16202 704960
rect 19954 703520 20066 704960
rect 23818 703520 23930 704960
rect 27682 703520 27794 704960
rect 31546 703520 31658 704960
rect 35410 703520 35522 704960
rect 39274 703520 39386 704960
rect 43138 703520 43250 704960
rect 47002 703520 47114 704960
rect 50866 703520 50978 704960
rect 54730 703520 54842 704960
rect 58594 703520 58706 704960
rect 62458 703520 62570 704960
rect 66322 703520 66434 704960
rect 70186 703520 70298 704960
rect 73406 703520 73518 704960
rect 77270 703520 77382 704960
rect 80072 703582 81020 703610
rect 12912 703474 12940 703520
rect 12728 703446 12940 703474
rect 16132 700398 16160 703520
rect 19996 700466 20024 703520
rect 23860 702434 23888 703520
rect 23492 702406 23888 702434
rect 19984 700460 20036 700466
rect 19984 700402 20036 700408
rect 16120 700392 16172 700398
rect 16120 700334 16172 700340
rect 14464 487212 14516 487218
rect 14464 487154 14516 487160
rect 14476 264314 14504 487154
rect 17224 483064 17276 483070
rect 17224 483006 17276 483012
rect 17236 271182 17264 483006
rect 17224 271176 17276 271182
rect 17224 271118 17276 271124
rect 14464 264308 14516 264314
rect 14464 264250 14516 264256
rect 23492 263498 23520 702406
rect 27724 683114 27752 703520
rect 31024 700460 31076 700466
rect 31024 700402 31076 700408
rect 27632 683086 27752 683114
rect 23480 263492 23532 263498
rect 23480 263434 23532 263440
rect 27632 193905 27660 683086
rect 31036 199481 31064 700402
rect 31588 700330 31616 703520
rect 35452 702434 35480 703520
rect 39316 702434 39344 703520
rect 43180 702434 43208 703520
rect 34532 702406 35480 702434
rect 38672 702406 39344 702434
rect 42812 702406 43208 702434
rect 31576 700324 31628 700330
rect 31576 700266 31628 700272
rect 31022 199472 31078 199481
rect 31022 199407 31078 199416
rect 27618 193896 27674 193905
rect 27618 193831 27674 193840
rect 34532 193225 34560 702406
rect 38672 265577 38700 702406
rect 38658 265568 38714 265577
rect 38658 265503 38714 265512
rect 34518 193216 34574 193225
rect 34518 193151 34574 193160
rect 12438 190224 12494 190233
rect 12438 190159 12494 190168
rect 42812 187649 42840 702406
rect 47044 683114 47072 703520
rect 50908 703050 50936 703520
rect 49700 703044 49752 703050
rect 49700 702986 49752 702992
rect 50896 703044 50948 703050
rect 50896 702986 50948 702992
rect 46952 683086 47072 683114
rect 46952 199510 46980 683086
rect 46940 199504 46992 199510
rect 46940 199446 46992 199452
rect 42798 187640 42854 187649
rect 42798 187575 42854 187584
rect 49712 186153 49740 702986
rect 54772 702434 54800 703520
rect 58636 702434 58664 703520
rect 62500 702434 62528 703520
rect 53852 702406 54800 702434
rect 57992 702406 58664 702434
rect 62132 702406 62528 702434
rect 53852 188358 53880 702406
rect 57992 263430 58020 702406
rect 61384 543788 61436 543794
rect 61384 543730 61436 543736
rect 57980 263424 58032 263430
rect 57980 263366 58032 263372
rect 61396 198014 61424 543730
rect 61384 198008 61436 198014
rect 61384 197950 61436 197956
rect 62132 197033 62160 702406
rect 66364 700534 66392 703520
rect 70228 703050 70256 703520
rect 69020 703044 69072 703050
rect 69020 702986 69072 702992
rect 70216 703044 70268 703050
rect 70216 702986 70268 702992
rect 66352 700528 66404 700534
rect 66352 700470 66404 700476
rect 69032 263362 69060 702986
rect 77312 700466 77340 703520
rect 78036 700528 78088 700534
rect 78036 700470 78088 700476
rect 77300 700460 77352 700466
rect 77300 700402 77352 700408
rect 77944 700392 77996 700398
rect 77944 700334 77996 700340
rect 75184 346452 75236 346458
rect 75184 346394 75236 346400
rect 75196 264382 75224 346394
rect 75184 264376 75236 264382
rect 75184 264318 75236 264324
rect 69020 263356 69072 263362
rect 69020 263298 69072 263304
rect 62118 197024 62174 197033
rect 62118 196959 62174 196968
rect 53840 188352 53892 188358
rect 77956 188329 77984 700334
rect 78048 200705 78076 700470
rect 78034 200696 78090 200705
rect 78034 200631 78090 200640
rect 80072 191214 80100 703582
rect 80992 703474 81020 703582
rect 81134 703520 81246 704960
rect 84212 703582 84884 703610
rect 81176 703474 81204 703520
rect 80992 703446 81204 703474
rect 80704 661088 80756 661094
rect 80704 661030 80756 661036
rect 80060 191208 80112 191214
rect 80060 191150 80112 191156
rect 53840 188294 53892 188300
rect 77942 188320 77998 188329
rect 77942 188255 77998 188264
rect 49698 186144 49754 186153
rect 49698 186079 49754 186088
rect 80716 183530 80744 661030
rect 84212 199578 84240 703582
rect 84856 703474 84884 703582
rect 84998 703520 85110 704960
rect 88862 703520 88974 704960
rect 92726 703520 92838 704960
rect 96590 703520 96702 704960
rect 100454 703520 100566 704960
rect 103532 703582 104204 703610
rect 85040 703474 85068 703520
rect 84856 703446 85068 703474
rect 92768 702434 92796 703520
rect 92492 702406 92796 702434
rect 88984 692844 89036 692850
rect 88984 692786 89036 692792
rect 84844 667956 84896 667962
rect 84844 667898 84896 667904
rect 84200 199572 84252 199578
rect 84200 199514 84252 199520
rect 84856 187610 84884 667898
rect 86224 600364 86276 600370
rect 86224 600306 86276 600312
rect 86236 192574 86264 600306
rect 86316 523048 86368 523054
rect 86316 522990 86368 522996
rect 86224 192568 86276 192574
rect 86224 192510 86276 192516
rect 84844 187604 84896 187610
rect 84844 187546 84896 187552
rect 80704 183524 80756 183530
rect 80704 183466 80756 183472
rect 86328 182850 86356 522990
rect 86408 443012 86460 443018
rect 86408 442954 86460 442960
rect 86420 185910 86448 442954
rect 88996 194041 89024 692786
rect 89076 688696 89128 688702
rect 89076 688638 89128 688644
rect 88982 194032 89038 194041
rect 88982 193967 89038 193976
rect 89088 191049 89116 688638
rect 90364 583772 90416 583778
rect 90364 583714 90416 583720
rect 89168 430636 89220 430642
rect 89168 430578 89220 430584
rect 89074 191040 89130 191049
rect 89074 190975 89130 190984
rect 89180 188426 89208 430578
rect 89260 378208 89312 378214
rect 89260 378150 89312 378156
rect 89168 188420 89220 188426
rect 89168 188362 89220 188368
rect 89272 185978 89300 378150
rect 90376 186182 90404 583714
rect 90456 571396 90508 571402
rect 90456 571338 90508 571344
rect 90468 193526 90496 571338
rect 91744 567248 91796 567254
rect 91744 567190 91796 567196
rect 90548 411324 90600 411330
rect 90548 411266 90600 411272
rect 90456 193520 90508 193526
rect 90456 193462 90508 193468
rect 90560 186998 90588 411266
rect 91756 190330 91784 567190
rect 91836 478916 91888 478922
rect 91836 478858 91888 478864
rect 91744 190324 91796 190330
rect 91744 190266 91796 190272
rect 91848 187678 91876 478858
rect 92492 202201 92520 702406
rect 94504 680400 94556 680406
rect 94504 680342 94556 680348
rect 93124 560312 93176 560318
rect 93124 560254 93176 560260
rect 92478 202192 92534 202201
rect 92478 202127 92534 202136
rect 93136 191690 93164 560254
rect 93216 495508 93268 495514
rect 93216 495450 93268 495456
rect 93124 191684 93176 191690
rect 93124 191626 93176 191632
rect 91836 187672 91888 187678
rect 91836 187614 91888 187620
rect 90548 186992 90600 186998
rect 90548 186934 90600 186940
rect 90364 186176 90416 186182
rect 90364 186118 90416 186124
rect 89260 185972 89312 185978
rect 89260 185914 89312 185920
rect 86408 185904 86460 185910
rect 86408 185846 86460 185852
rect 93228 185842 93256 495450
rect 93308 407176 93360 407182
rect 93308 407118 93360 407124
rect 93320 192642 93348 407118
rect 93308 192636 93360 192642
rect 93308 192578 93360 192584
rect 94516 188873 94544 680342
rect 95884 627972 95936 627978
rect 95884 627914 95936 627920
rect 94596 531344 94648 531350
rect 94596 531286 94648 531292
rect 94608 194274 94636 531286
rect 94688 455456 94740 455462
rect 94688 455398 94740 455404
rect 94596 194268 94648 194274
rect 94596 194210 94648 194216
rect 94596 193928 94648 193934
rect 94596 193870 94648 193876
rect 94502 188864 94558 188873
rect 94502 188799 94558 188808
rect 93216 185836 93268 185842
rect 93216 185778 93268 185784
rect 86316 182844 86368 182850
rect 86316 182786 86368 182792
rect 82820 142860 82872 142866
rect 82820 142802 82872 142808
rect 59360 142384 59412 142390
rect 59360 142326 59412 142332
rect 3516 141364 3568 141370
rect 3516 141306 3568 141312
rect 8944 141364 8996 141370
rect 8944 141306 8996 141312
rect 3528 140865 3556 141306
rect 3514 140856 3570 140865
rect 3514 140791 3570 140800
rect 4804 140820 4856 140826
rect 4804 140762 4856 140768
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136678 3464 136711
rect 3424 136672 3476 136678
rect 3424 136614 3476 136620
rect 3148 121440 3200 121446
rect 3148 121382 3200 121388
rect 3160 120465 3188 121382
rect 3146 120456 3202 120465
rect 3146 120391 3202 120400
rect 3240 117292 3292 117298
rect 3240 117234 3292 117240
rect 3252 117065 3280 117234
rect 3238 117056 3294 117065
rect 3238 116991 3294 117000
rect 3422 112976 3478 112985
rect 3422 112911 3478 112920
rect 3436 111858 3464 112911
rect 3424 111852 3476 111858
rect 3424 111794 3476 111800
rect 3424 108996 3476 109002
rect 3424 108938 3476 108944
rect 3436 108905 3464 108938
rect 3422 108896 3478 108905
rect 3422 108831 3478 108840
rect 3422 104816 3478 104825
rect 3422 104751 3478 104760
rect 3436 103562 3464 104751
rect 3424 103556 3476 103562
rect 3424 103498 3476 103504
rect 3330 100736 3386 100745
rect 3330 100671 3386 100680
rect 3344 93854 3372 100671
rect 3424 96688 3476 96694
rect 3422 96656 3424 96665
rect 3476 96656 3478 96665
rect 3422 96591 3478 96600
rect 3148 93832 3200 93838
rect 3344 93826 3556 93854
rect 3148 93774 3200 93780
rect 3160 92585 3188 93774
rect 3146 92576 3202 92585
rect 3146 92511 3202 92520
rect 3422 84416 3478 84425
rect 3422 84351 3478 84360
rect 3436 84250 3464 84351
rect 3424 84244 3476 84250
rect 3424 84186 3476 84192
rect 3424 81388 3476 81394
rect 3424 81330 3476 81336
rect 3436 80345 3464 81330
rect 3422 80336 3478 80345
rect 3422 80271 3478 80280
rect 3528 79354 3556 93826
rect 3516 79348 3568 79354
rect 3516 79290 3568 79296
rect 4816 77246 4844 140762
rect 2780 77240 2832 77246
rect 2780 77182 2832 77188
rect 4804 77240 4856 77246
rect 4804 77182 4856 77188
rect 2792 76265 2820 77182
rect 2778 76256 2834 76265
rect 2778 76191 2834 76200
rect 36544 75268 36596 75274
rect 36544 75210 36596 75216
rect 13084 73840 13136 73846
rect 13084 73782 13136 73788
rect 3148 73160 3200 73166
rect 3148 73102 3200 73108
rect 3160 72185 3188 73102
rect 3146 72176 3202 72185
rect 3146 72111 3202 72120
rect 4804 71052 4856 71058
rect 4804 70994 4856 71000
rect 3148 68944 3200 68950
rect 3148 68886 3200 68892
rect 3160 68105 3188 68886
rect 3146 68096 3202 68105
rect 3146 68031 3202 68040
rect 3148 64864 3200 64870
rect 3148 64806 3200 64812
rect 3160 64025 3188 64806
rect 3146 64016 3202 64025
rect 3146 63951 3202 63960
rect 3424 56568 3476 56574
rect 3422 56536 3424 56545
rect 3476 56536 3478 56545
rect 3422 56471 3478 56480
rect 3516 53100 3568 53106
rect 3516 53042 3568 53048
rect 3422 52456 3478 52465
rect 3422 52391 3424 52400
rect 3476 52391 3478 52400
rect 3424 52362 3476 52368
rect 3240 49700 3292 49706
rect 3240 49642 3292 49648
rect 3252 48385 3280 49642
rect 3528 49314 3556 53042
rect 3436 49286 3556 49314
rect 3238 48376 3294 48385
rect 3238 48311 3294 48320
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 3160 36145 3188 37198
rect 3146 36136 3202 36145
rect 3146 36071 3202 36080
rect 3148 33040 3200 33046
rect 3148 32982 3200 32988
rect 3160 32065 3188 32982
rect 3146 32056 3202 32065
rect 3146 31991 3202 32000
rect 3148 28960 3200 28966
rect 3148 28902 3200 28908
rect 3160 27985 3188 28902
rect 3146 27976 3202 27985
rect 3146 27911 3202 27920
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 3068 23905 3096 24754
rect 3054 23896 3110 23905
rect 3054 23831 3110 23840
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3068 11665 3096 12378
rect 3054 11656 3110 11665
rect 3054 11591 3110 11600
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7585 3004 8230
rect 2962 7576 3018 7585
rect 2962 7511 3018 7520
rect 3436 6914 3464 49286
rect 3516 45552 3568 45558
rect 3516 45494 3568 45500
rect 3528 44305 3556 45494
rect 3514 44296 3570 44305
rect 3514 44231 3570 44240
rect 3516 41404 3568 41410
rect 3516 41346 3568 41352
rect 3528 40225 3556 41346
rect 3514 40216 3570 40225
rect 3514 40151 3570 40160
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19825 3556 20606
rect 3514 19816 3570 19825
rect 3514 19751 3570 19760
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15745 3556 16526
rect 3514 15736 3570 15745
rect 3514 15671 3570 15680
rect 3344 6886 3464 6914
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 20 3596 72 3602
rect 20 3538 72 3544
rect 32 480 60 3538
rect 3160 3505 3188 4082
rect 3344 3602 3372 6886
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 4816 3534 4844 70994
rect 6920 57248 6972 57254
rect 6920 57190 6972 57196
rect 6932 16574 6960 57190
rect 6932 16546 7144 16574
rect 3240 3528 3292 3534
rect 3146 3496 3202 3505
rect 3240 3470 3292 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3146 3431 3202 3440
rect 3252 480 3280 3470
rect 7116 480 7144 16546
rect 13096 8294 13124 73782
rect 26240 66904 26292 66910
rect 26240 66846 26292 66852
rect 22744 61396 22796 61402
rect 22744 61338 22796 61344
rect 17960 55956 18012 55962
rect 17960 55898 18012 55904
rect 13820 54528 13872 54534
rect 13820 54470 13872 54476
rect 13832 16574 13860 54470
rect 17972 16574 18000 55898
rect 22756 45558 22784 61338
rect 22744 45552 22796 45558
rect 22744 45494 22796 45500
rect 26252 16574 26280 66846
rect 35164 65544 35216 65550
rect 35164 65486 35216 65492
rect 31024 62892 31076 62898
rect 31024 62834 31076 62840
rect 13832 16546 14872 16574
rect 17972 16546 18736 16574
rect 26252 16546 26464 16574
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 14844 480 14872 16546
rect 18708 480 18736 16546
rect 26436 480 26464 16546
rect 31036 3534 31064 62834
rect 35176 24818 35204 65486
rect 35164 24812 35216 24818
rect 35164 24754 35216 24760
rect 36556 3738 36584 75210
rect 54484 72480 54536 72486
rect 54484 72422 54536 72428
rect 43444 69692 43496 69698
rect 43444 69634 43496 69640
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 34152 3732 34204 3738
rect 34152 3674 34204 3680
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 30300 480 30328 3470
rect 34164 480 34192 3674
rect 38028 480 38056 4762
rect 43456 3534 43484 69634
rect 48320 60036 48372 60042
rect 48320 59978 48372 59984
rect 48332 3534 48360 59978
rect 54496 4146 54524 72422
rect 59372 16574 59400 142326
rect 67640 76560 67692 76566
rect 67640 76502 67692 76508
rect 64144 69760 64196 69766
rect 64144 69702 64196 69708
rect 59372 16546 60136 16574
rect 54484 4140 54536 4146
rect 54484 4082 54536 4088
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 48320 3528 48372 3534
rect 48320 3470 48372 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 53472 3528 53524 3534
rect 53472 3470 53524 3476
rect 41892 480 41920 3470
rect 49620 480 49648 3470
rect 53484 480 53512 3470
rect -10 -960 102 480
rect 3210 -960 3322 480
rect 7074 -960 7186 480
rect 10938 -960 11050 480
rect 14802 -960 14914 480
rect 18666 -960 18778 480
rect 22530 -960 22642 480
rect 26394 -960 26506 480
rect 30258 -960 30370 480
rect 34122 -960 34234 480
rect 37986 -960 38098 480
rect 41850 -960 41962 480
rect 45714 -960 45826 480
rect 49578 -960 49690 480
rect 53442 -960 53554 480
rect 56662 -960 56774 480
rect 60108 354 60136 16546
rect 64156 3534 64184 69702
rect 67652 16574 67680 76502
rect 78680 75200 78732 75206
rect 78680 75142 78732 75148
rect 78692 16574 78720 75142
rect 82832 16574 82860 142802
rect 94608 72282 94636 193870
rect 94700 191282 94728 455398
rect 94780 321632 94832 321638
rect 94780 321574 94832 321580
rect 94688 191276 94740 191282
rect 94688 191218 94740 191224
rect 94792 188834 94820 321574
rect 94872 317484 94924 317490
rect 94872 317426 94924 317432
rect 94780 188828 94832 188834
rect 94780 188770 94832 188776
rect 94884 188766 94912 317426
rect 95148 200864 95200 200870
rect 95148 200806 95200 200812
rect 95054 200696 95110 200705
rect 95054 200631 95110 200640
rect 94964 200320 95016 200326
rect 94964 200262 95016 200268
rect 94872 188760 94924 188766
rect 94872 188702 94924 188708
rect 94780 181484 94832 181490
rect 94780 181426 94832 181432
rect 94792 180878 94820 181426
rect 94780 180872 94832 180878
rect 94780 180814 94832 180820
rect 94688 172576 94740 172582
rect 94688 172518 94740 172524
rect 94700 76362 94728 172518
rect 94688 76356 94740 76362
rect 94688 76298 94740 76304
rect 94792 73710 94820 180814
rect 94872 173188 94924 173194
rect 94872 173130 94924 173136
rect 94884 172582 94912 173130
rect 94872 172576 94924 172582
rect 94872 172518 94924 172524
rect 94976 76634 95004 200262
rect 95068 200161 95096 200631
rect 95160 200190 95188 200806
rect 95148 200184 95200 200190
rect 95054 200152 95110 200161
rect 95148 200126 95200 200132
rect 95054 200087 95110 200096
rect 94964 76628 95016 76634
rect 94964 76570 95016 76576
rect 94780 73704 94832 73710
rect 94780 73646 94832 73652
rect 94596 72276 94648 72282
rect 94596 72218 94648 72224
rect 95068 68882 95096 200087
rect 95056 68876 95108 68882
rect 95056 68818 95108 68824
rect 95160 65346 95188 200126
rect 95896 188494 95924 627914
rect 95976 587920 96028 587926
rect 95976 587862 96028 587868
rect 95884 188488 95936 188494
rect 95884 188430 95936 188436
rect 95988 184686 96016 587862
rect 96344 512032 96396 512038
rect 96344 511974 96396 511980
rect 96160 403028 96212 403034
rect 96160 402970 96212 402976
rect 96068 201544 96120 201550
rect 96068 201486 96120 201492
rect 95976 184680 96028 184686
rect 95976 184622 96028 184628
rect 95976 141568 96028 141574
rect 95976 141510 96028 141516
rect 95988 74534 96016 141510
rect 96080 79490 96108 201486
rect 96172 183394 96200 402970
rect 96252 200864 96304 200870
rect 96252 200806 96304 200812
rect 96160 183388 96212 183394
rect 96160 183330 96212 183336
rect 96068 79484 96120 79490
rect 96068 79426 96120 79432
rect 95988 74506 96108 74534
rect 95148 65340 95200 65346
rect 95148 65282 95200 65288
rect 96080 60722 96108 74506
rect 96172 63510 96200 183330
rect 96264 77790 96292 200806
rect 96356 195265 96384 511974
rect 96436 200796 96488 200802
rect 96436 200738 96488 200744
rect 96448 200258 96476 200738
rect 96436 200252 96488 200258
rect 96436 200194 96488 200200
rect 96342 195256 96398 195265
rect 96342 195191 96398 195200
rect 96344 194608 96396 194614
rect 96344 194550 96396 194556
rect 96252 77784 96304 77790
rect 96252 77726 96304 77732
rect 96356 64802 96384 194550
rect 96448 67590 96476 200194
rect 96528 196716 96580 196722
rect 96528 196658 96580 196664
rect 96436 67584 96488 67590
rect 96436 67526 96488 67532
rect 96344 64796 96396 64802
rect 96344 64738 96396 64744
rect 96160 63504 96212 63510
rect 96160 63446 96212 63452
rect 96540 63306 96568 196658
rect 96632 193322 96660 703520
rect 98644 701072 98696 701078
rect 98644 701014 98696 701020
rect 97264 612808 97316 612814
rect 97264 612750 97316 612756
rect 96620 193316 96672 193322
rect 96620 193258 96672 193264
rect 96632 190454 96660 193258
rect 97276 191486 97304 612750
rect 97356 499588 97408 499594
rect 97356 499530 97408 499536
rect 97368 197266 97396 499530
rect 97448 361616 97500 361622
rect 97448 361558 97500 361564
rect 97356 197260 97408 197266
rect 97356 197202 97408 197208
rect 97460 191554 97488 361558
rect 97816 277432 97868 277438
rect 97816 277374 97868 277380
rect 97540 200388 97592 200394
rect 97540 200330 97592 200336
rect 97448 191548 97500 191554
rect 97448 191490 97500 191496
rect 97264 191480 97316 191486
rect 97264 191422 97316 191428
rect 96632 190426 97028 190454
rect 97000 75041 97028 190426
rect 97356 189712 97408 189718
rect 97356 189654 97408 189660
rect 97264 142996 97316 143002
rect 97264 142938 97316 142944
rect 97078 141808 97134 141817
rect 97078 141743 97134 141752
rect 97092 75721 97120 141743
rect 97172 140072 97224 140078
rect 97172 140014 97224 140020
rect 97078 75712 97134 75721
rect 97078 75647 97134 75656
rect 96986 75032 97042 75041
rect 96986 74967 97042 74976
rect 97184 63442 97212 140014
rect 97172 63436 97224 63442
rect 97172 63378 97224 63384
rect 96528 63300 96580 63306
rect 96528 63242 96580 63248
rect 96068 60716 96120 60722
rect 96068 60658 96120 60664
rect 93124 60104 93176 60110
rect 93124 60046 93176 60052
rect 67652 16546 67864 16574
rect 78692 16546 79456 16574
rect 82832 16546 83320 16574
rect 64144 3528 64196 3534
rect 64144 3470 64196 3476
rect 64420 3460 64472 3466
rect 64420 3402 64472 3408
rect 64432 480 64460 3402
rect 60526 354 60638 480
rect 60108 326 60638 354
rect 60526 -960 60638 326
rect 64390 -960 64502 480
rect 67836 354 67864 16546
rect 72148 3528 72200 3534
rect 72148 3470 72200 3476
rect 72160 480 72188 3470
rect 68254 354 68366 480
rect 67836 326 68366 354
rect 68254 -960 68366 326
rect 72118 -960 72230 480
rect 75982 -960 76094 480
rect 79428 354 79456 16546
rect 79846 354 79958 480
rect 79428 326 79958 354
rect 83292 354 83320 16546
rect 93136 3602 93164 60046
rect 96080 60042 96108 60658
rect 96068 60036 96120 60042
rect 96068 59978 96120 59984
rect 95240 58676 95292 58682
rect 95240 58618 95292 58624
rect 95252 16574 95280 58618
rect 97276 56574 97304 142938
rect 97368 75818 97396 189654
rect 97552 79694 97580 200330
rect 97724 198552 97776 198558
rect 97724 198494 97776 198500
rect 97630 191176 97686 191185
rect 97630 191111 97686 191120
rect 97540 79688 97592 79694
rect 97540 79630 97592 79636
rect 97356 75812 97408 75818
rect 97356 75754 97408 75760
rect 97644 64841 97672 191111
rect 97736 67561 97764 198494
rect 97828 186046 97856 277374
rect 98656 193089 98684 701014
rect 98736 644496 98788 644502
rect 98736 644438 98788 644444
rect 98642 193080 98698 193089
rect 98642 193015 98698 193024
rect 98748 188698 98776 644438
rect 98828 615528 98880 615534
rect 98828 615470 98880 615476
rect 98736 188692 98788 188698
rect 98736 188634 98788 188640
rect 98840 188601 98868 615470
rect 102784 604512 102836 604518
rect 102784 604454 102836 604460
rect 101404 596216 101456 596222
rect 101404 596158 101456 596164
rect 100024 579692 100076 579698
rect 100024 579634 100076 579640
rect 98920 422340 98972 422346
rect 98920 422282 98972 422288
rect 98826 188592 98882 188601
rect 98826 188527 98882 188536
rect 97816 186040 97868 186046
rect 97816 185982 97868 185988
rect 98828 185632 98880 185638
rect 98828 185574 98880 185580
rect 98644 151156 98696 151162
rect 98644 151098 98696 151104
rect 97908 148368 97960 148374
rect 97908 148310 97960 148316
rect 97816 143608 97868 143614
rect 97816 143550 97868 143556
rect 97722 67552 97778 67561
rect 97722 67487 97778 67496
rect 97630 64832 97686 64841
rect 97630 64767 97686 64776
rect 97264 56568 97316 56574
rect 97264 56510 97316 56516
rect 95252 16546 95372 16574
rect 91468 3596 91520 3602
rect 91468 3538 91520 3544
rect 93124 3596 93176 3602
rect 93124 3538 93176 3544
rect 91480 480 91508 3538
rect 95344 480 95372 16546
rect 97828 3602 97856 143550
rect 97920 69018 97948 148310
rect 98000 143268 98052 143274
rect 98000 143210 98052 143216
rect 97908 69012 97960 69018
rect 97908 68954 97960 68960
rect 98012 16574 98040 143210
rect 98552 84244 98604 84250
rect 98552 84186 98604 84192
rect 98564 71097 98592 84186
rect 98656 72418 98684 151098
rect 98736 148640 98788 148646
rect 98736 148582 98788 148588
rect 98644 72412 98696 72418
rect 98644 72354 98696 72360
rect 98550 71088 98606 71097
rect 98550 71023 98606 71032
rect 98748 69766 98776 148582
rect 98840 78878 98868 185574
rect 98932 184754 98960 422282
rect 99932 273284 99984 273290
rect 99932 273226 99984 273232
rect 99288 198008 99340 198014
rect 99288 197950 99340 197956
rect 99012 192568 99064 192574
rect 99012 192510 99064 192516
rect 98920 184748 98972 184754
rect 98920 184690 98972 184696
rect 98920 177404 98972 177410
rect 98920 177346 98972 177352
rect 98828 78872 98880 78878
rect 98828 78814 98880 78820
rect 98736 69760 98788 69766
rect 98736 69702 98788 69708
rect 98932 67289 98960 177346
rect 99024 81161 99052 192510
rect 99104 191140 99156 191146
rect 99104 191082 99156 191088
rect 99010 81152 99066 81161
rect 99010 81087 99066 81096
rect 99116 77586 99144 191082
rect 99194 188320 99250 188329
rect 99194 188255 99250 188264
rect 99104 77580 99156 77586
rect 99104 77522 99156 77528
rect 99208 74225 99236 188255
rect 99194 74216 99250 74225
rect 99194 74151 99250 74160
rect 99300 69562 99328 197950
rect 99944 184550 99972 273226
rect 100036 188902 100064 579634
rect 100116 459604 100168 459610
rect 100116 459546 100168 459552
rect 100128 191350 100156 459546
rect 100208 386436 100260 386442
rect 100208 386378 100260 386384
rect 100220 191826 100248 386378
rect 100300 354748 100352 354754
rect 100300 354690 100352 354696
rect 100208 191820 100260 191826
rect 100208 191762 100260 191768
rect 100208 191412 100260 191418
rect 100208 191354 100260 191360
rect 100116 191344 100168 191350
rect 100116 191286 100168 191292
rect 100220 190534 100248 191354
rect 100208 190528 100260 190534
rect 100208 190470 100260 190476
rect 100024 188896 100076 188902
rect 100024 188838 100076 188844
rect 99932 184544 99984 184550
rect 99932 184486 99984 184492
rect 100116 176724 100168 176730
rect 100116 176666 100168 176672
rect 99932 151292 99984 151298
rect 99932 151234 99984 151240
rect 99840 151088 99892 151094
rect 99840 151030 99892 151036
rect 99288 69556 99340 69562
rect 99288 69498 99340 69504
rect 98918 67280 98974 67289
rect 98918 67215 98974 67224
rect 99852 65482 99880 151030
rect 99944 65822 99972 151234
rect 100024 151224 100076 151230
rect 100024 151166 100076 151172
rect 100036 65958 100064 151166
rect 100128 69873 100156 176666
rect 100220 81977 100248 190470
rect 100312 188630 100340 354690
rect 100668 198348 100720 198354
rect 100668 198290 100720 198296
rect 100392 198212 100444 198218
rect 100392 198154 100444 198160
rect 100300 188624 100352 188630
rect 100300 188566 100352 188572
rect 100300 187060 100352 187066
rect 100300 187002 100352 187008
rect 100206 81968 100262 81977
rect 100206 81903 100262 81912
rect 100312 72486 100340 187002
rect 100404 75886 100432 198154
rect 100576 198076 100628 198082
rect 100576 198018 100628 198024
rect 100484 195424 100536 195430
rect 100484 195366 100536 195372
rect 100392 75880 100444 75886
rect 100392 75822 100444 75828
rect 100300 72480 100352 72486
rect 100300 72422 100352 72428
rect 100114 69864 100170 69873
rect 100114 69799 100170 69808
rect 100024 65952 100076 65958
rect 100024 65894 100076 65900
rect 99932 65816 99984 65822
rect 99932 65758 99984 65764
rect 99840 65476 99892 65482
rect 99840 65418 99892 65424
rect 100496 63374 100524 195366
rect 100588 64666 100616 198018
rect 100576 64660 100628 64666
rect 100576 64602 100628 64608
rect 100680 64530 100708 198290
rect 101416 183462 101444 596158
rect 101496 294024 101548 294030
rect 101496 293966 101548 293972
rect 101508 184618 101536 293966
rect 102692 281580 102744 281586
rect 102692 281522 102744 281528
rect 102048 198416 102100 198422
rect 102048 198358 102100 198364
rect 101956 198280 102008 198286
rect 101956 198222 102008 198228
rect 101864 192636 101916 192642
rect 101864 192578 101916 192584
rect 101772 191888 101824 191894
rect 101772 191830 101824 191836
rect 101496 184612 101548 184618
rect 101496 184554 101548 184560
rect 101404 183456 101456 183462
rect 101404 183398 101456 183404
rect 101588 177472 101640 177478
rect 101588 177414 101640 177420
rect 101496 177336 101548 177342
rect 101496 177278 101548 177284
rect 101220 148708 101272 148714
rect 101220 148650 101272 148656
rect 101232 79762 101260 148650
rect 101404 148504 101456 148510
rect 101404 148446 101456 148452
rect 101312 147008 101364 147014
rect 101312 146950 101364 146956
rect 101220 79756 101272 79762
rect 101220 79698 101272 79704
rect 101324 65890 101352 146950
rect 101312 65884 101364 65890
rect 101312 65826 101364 65832
rect 100668 64524 100720 64530
rect 100668 64466 100720 64472
rect 100484 63368 100536 63374
rect 100484 63310 100536 63316
rect 101416 55214 101444 148446
rect 101508 81025 101536 177278
rect 101494 81016 101550 81025
rect 101494 80951 101550 80960
rect 101600 79121 101628 177414
rect 101680 175976 101732 175982
rect 101680 175918 101732 175924
rect 101586 79112 101642 79121
rect 101586 79047 101642 79056
rect 101692 77217 101720 175918
rect 101678 77208 101734 77217
rect 101678 77143 101734 77152
rect 101784 70922 101812 191830
rect 101772 70916 101824 70922
rect 101772 70858 101824 70864
rect 101876 68610 101904 192578
rect 101968 72894 101996 198222
rect 101956 72888 102008 72894
rect 101956 72830 102008 72836
rect 101864 68604 101916 68610
rect 101864 68546 101916 68552
rect 102060 65686 102088 198358
rect 102600 193996 102652 194002
rect 102600 193938 102652 193944
rect 102612 109002 102640 193938
rect 102704 191622 102732 281522
rect 102692 191616 102744 191622
rect 102692 191558 102744 191564
rect 102796 188154 102824 604454
rect 102876 575544 102928 575550
rect 102876 575486 102928 575492
rect 102784 188148 102836 188154
rect 102784 188090 102836 188096
rect 102888 186318 102916 575486
rect 102968 516180 103020 516186
rect 102968 516122 103020 516128
rect 102980 195809 103008 516122
rect 103060 426488 103112 426494
rect 103060 426430 103112 426436
rect 102966 195800 103022 195809
rect 102966 195735 103022 195744
rect 103072 194206 103100 426430
rect 103152 419552 103204 419558
rect 103152 419494 103204 419500
rect 103164 194342 103192 419494
rect 103428 198484 103480 198490
rect 103428 198426 103480 198432
rect 103152 194336 103204 194342
rect 103152 194278 103204 194284
rect 103060 194200 103112 194206
rect 103060 194142 103112 194148
rect 103336 192704 103388 192710
rect 103336 192646 103388 192652
rect 103244 191752 103296 191758
rect 103244 191694 103296 191700
rect 102876 186312 102928 186318
rect 102876 186254 102928 186260
rect 103152 181620 103204 181626
rect 103152 181562 103204 181568
rect 103060 180872 103112 180878
rect 103060 180814 103112 180820
rect 102968 180192 103020 180198
rect 102968 180134 103020 180140
rect 102876 180124 102928 180130
rect 102876 180066 102928 180072
rect 102692 146940 102744 146946
rect 102692 146882 102744 146888
rect 102140 108996 102192 109002
rect 102140 108938 102192 108944
rect 102600 108996 102652 109002
rect 102600 108938 102652 108944
rect 102152 108322 102180 108938
rect 102140 108316 102192 108322
rect 102140 108258 102192 108264
rect 102704 81841 102732 146882
rect 102784 140344 102836 140350
rect 102784 140286 102836 140292
rect 102690 81832 102746 81841
rect 102690 81767 102746 81776
rect 102140 76492 102192 76498
rect 102140 76434 102192 76440
rect 102152 75886 102180 76434
rect 102140 75880 102192 75886
rect 102140 75822 102192 75828
rect 102048 65680 102100 65686
rect 102048 65622 102100 65628
rect 101404 55208 101456 55214
rect 101404 55150 101456 55156
rect 101416 54534 101444 55150
rect 101404 54528 101456 54534
rect 101404 54470 101456 54476
rect 102152 16574 102180 75822
rect 102796 66162 102824 140286
rect 102888 78985 102916 180066
rect 102980 79529 103008 180134
rect 102966 79520 103022 79529
rect 102966 79455 103022 79464
rect 102874 78976 102930 78985
rect 102874 78911 102930 78920
rect 103072 68134 103100 180814
rect 103060 68128 103112 68134
rect 103060 68070 103112 68076
rect 103164 66910 103192 181562
rect 103256 75546 103284 191694
rect 103244 75540 103296 75546
rect 103244 75482 103296 75488
rect 103152 66904 103204 66910
rect 103152 66846 103204 66852
rect 102784 66156 102836 66162
rect 102784 66098 102836 66104
rect 103348 64569 103376 192646
rect 103440 66842 103468 198426
rect 103532 193934 103560 703582
rect 104176 703474 104204 703582
rect 104318 703520 104430 704960
rect 107672 703582 108068 703610
rect 104360 703474 104388 703520
rect 104176 703446 104388 703474
rect 105544 672104 105596 672110
rect 105544 672046 105596 672052
rect 104164 539640 104216 539646
rect 104164 539582 104216 539588
rect 103612 451308 103664 451314
rect 103612 451250 103664 451256
rect 103624 194614 103652 451250
rect 103612 194608 103664 194614
rect 103612 194550 103664 194556
rect 103520 193928 103572 193934
rect 103520 193870 103572 193876
rect 104176 193254 104204 539582
rect 104256 350600 104308 350606
rect 104256 350542 104308 350548
rect 104268 197062 104296 350542
rect 104900 342304 104952 342310
rect 104900 342246 104952 342252
rect 104532 200524 104584 200530
rect 104532 200466 104584 200472
rect 104440 200456 104492 200462
rect 104440 200398 104492 200404
rect 104256 197056 104308 197062
rect 104256 196998 104308 197004
rect 104348 194540 104400 194546
rect 104348 194482 104400 194488
rect 104360 193934 104388 194482
rect 104348 193928 104400 193934
rect 104348 193870 104400 193876
rect 104164 193248 104216 193254
rect 104164 193190 104216 193196
rect 104348 186312 104400 186318
rect 104348 186254 104400 186260
rect 104360 185706 104388 186254
rect 104348 185700 104400 185706
rect 104348 185642 104400 185648
rect 104360 184226 104388 185642
rect 104176 184198 104388 184226
rect 104072 148844 104124 148850
rect 104072 148786 104124 148792
rect 103980 140140 104032 140146
rect 103980 140082 104032 140088
rect 103992 117298 104020 140082
rect 103980 117292 104032 117298
rect 103980 117234 104032 117240
rect 103992 77994 104020 117234
rect 104084 78470 104112 148786
rect 104072 78464 104124 78470
rect 104072 78406 104124 78412
rect 103980 77988 104032 77994
rect 103980 77930 104032 77936
rect 104176 72729 104204 184198
rect 104348 184136 104400 184142
rect 104348 184078 104400 184084
rect 104256 181688 104308 181694
rect 104256 181630 104308 181636
rect 104162 72720 104218 72729
rect 104162 72655 104218 72664
rect 103428 66836 103480 66842
rect 103428 66778 103480 66784
rect 103334 64560 103390 64569
rect 103334 64495 103390 64504
rect 104268 64462 104296 181630
rect 104360 67046 104388 184078
rect 104452 78402 104480 200398
rect 104544 78538 104572 200466
rect 104808 196920 104860 196926
rect 104808 196862 104860 196868
rect 104714 195392 104770 195401
rect 104714 195327 104770 195336
rect 104624 194608 104676 194614
rect 104624 194550 104676 194556
rect 104636 194138 104664 194550
rect 104624 194132 104676 194138
rect 104624 194074 104676 194080
rect 104624 193928 104676 193934
rect 104624 193870 104676 193876
rect 104532 78532 104584 78538
rect 104532 78474 104584 78480
rect 104440 78396 104492 78402
rect 104440 78338 104492 78344
rect 104636 67386 104664 193870
rect 104624 67380 104676 67386
rect 104624 67322 104676 67328
rect 104728 67318 104756 195327
rect 104820 68746 104848 196862
rect 104912 189718 104940 342246
rect 105556 196897 105584 672046
rect 106924 619676 106976 619682
rect 106924 619618 106976 619624
rect 105636 358828 105688 358834
rect 105636 358770 105688 358776
rect 105648 200297 105676 358770
rect 105728 305040 105780 305046
rect 105728 304982 105780 304988
rect 105634 200288 105690 200297
rect 105634 200223 105690 200232
rect 105542 196888 105598 196897
rect 105542 196823 105598 196832
rect 105648 191894 105676 200223
rect 105740 194954 105768 304982
rect 106832 264988 106884 264994
rect 106832 264930 106884 264936
rect 106188 198144 106240 198150
rect 106188 198086 106240 198092
rect 105728 194948 105780 194954
rect 105728 194890 105780 194896
rect 105636 191888 105688 191894
rect 105636 191830 105688 191836
rect 104900 189712 104952 189718
rect 104900 189654 104952 189660
rect 105820 189236 105872 189242
rect 105820 189178 105872 189184
rect 105636 187808 105688 187814
rect 105636 187750 105688 187756
rect 105544 178696 105596 178702
rect 105544 178638 105596 178644
rect 105452 141908 105504 141914
rect 105452 141850 105504 141856
rect 105360 136672 105412 136678
rect 105360 136614 105412 136620
rect 104808 68740 104860 68746
rect 104808 68682 104860 68688
rect 104716 67312 104768 67318
rect 104716 67254 104768 67260
rect 104348 67040 104400 67046
rect 104348 66982 104400 66988
rect 105372 65754 105400 136614
rect 105360 65748 105412 65754
rect 105360 65690 105412 65696
rect 104256 64456 104308 64462
rect 104256 64398 104308 64404
rect 105464 53786 105492 141850
rect 105556 73574 105584 178638
rect 105648 80850 105676 187750
rect 105728 178764 105780 178770
rect 105728 178706 105780 178712
rect 105636 80844 105688 80850
rect 105636 80786 105688 80792
rect 105544 73568 105596 73574
rect 105544 73510 105596 73516
rect 105740 70961 105768 178706
rect 105832 79257 105860 189178
rect 105912 184408 105964 184414
rect 105912 184350 105964 184356
rect 105818 79248 105874 79257
rect 105818 79183 105874 79192
rect 105726 70952 105782 70961
rect 105726 70887 105782 70896
rect 105924 68678 105952 184350
rect 106096 184000 106148 184006
rect 106096 183942 106148 183948
rect 106004 181756 106056 181762
rect 106004 181698 106056 181704
rect 105912 68672 105964 68678
rect 105912 68614 105964 68620
rect 106016 64258 106044 181698
rect 106108 66706 106136 183942
rect 106096 66700 106148 66706
rect 106096 66642 106148 66648
rect 106200 64598 106228 198086
rect 106844 185570 106872 264930
rect 106936 191729 106964 619618
rect 107016 547936 107068 547942
rect 107016 547878 107068 547884
rect 107028 194478 107056 547878
rect 107200 472048 107252 472054
rect 107200 471990 107252 471996
rect 107108 463752 107160 463758
rect 107108 463694 107160 463700
rect 107016 194472 107068 194478
rect 107016 194414 107068 194420
rect 106922 191720 106978 191729
rect 106922 191655 106978 191664
rect 107120 191010 107148 463694
rect 107212 209774 107240 471990
rect 107212 209746 107608 209774
rect 107382 202192 107438 202201
rect 107382 202127 107438 202136
rect 107396 201521 107424 202127
rect 107382 201512 107438 201521
rect 107382 201447 107438 201456
rect 107292 197056 107344 197062
rect 107292 196998 107344 197004
rect 107108 191004 107160 191010
rect 107108 190946 107160 190952
rect 107200 188352 107252 188358
rect 107200 188294 107252 188300
rect 107212 187542 107240 188294
rect 107200 187536 107252 187542
rect 107200 187478 107252 187484
rect 106832 185564 106884 185570
rect 106832 185506 106884 185512
rect 107108 182232 107160 182238
rect 107108 182174 107160 182180
rect 106924 148980 106976 148986
rect 106924 148922 106976 148928
rect 106832 148912 106884 148918
rect 106832 148854 106884 148860
rect 106740 141432 106792 141438
rect 106740 141374 106792 141380
rect 106752 121446 106780 141374
rect 106740 121440 106792 121446
rect 106740 121382 106792 121388
rect 106844 78334 106872 148854
rect 106832 78328 106884 78334
rect 106832 78270 106884 78276
rect 106936 78130 106964 148922
rect 107016 148436 107068 148442
rect 107016 148378 107068 148384
rect 106924 78124 106976 78130
rect 106924 78066 106976 78072
rect 106280 72888 106332 72894
rect 106280 72830 106332 72836
rect 106188 64592 106240 64598
rect 106188 64534 106240 64540
rect 106004 64252 106056 64258
rect 106004 64194 106056 64200
rect 105452 53780 105504 53786
rect 105452 53722 105504 53728
rect 105464 53106 105492 53722
rect 105452 53100 105504 53106
rect 105452 53042 105504 53048
rect 106292 16574 106320 72830
rect 107028 68542 107056 148378
rect 107016 68536 107068 68542
rect 107016 68478 107068 68484
rect 107120 68377 107148 182174
rect 107212 68406 107240 187478
rect 107304 74526 107332 196998
rect 107396 190454 107424 201447
rect 107580 199306 107608 209746
rect 107568 199300 107620 199306
rect 107568 199242 107620 199248
rect 107396 190426 107516 190454
rect 107384 189780 107436 189786
rect 107384 189722 107436 189728
rect 107292 74520 107344 74526
rect 107292 74462 107344 74468
rect 107200 68400 107252 68406
rect 107106 68368 107162 68377
rect 107200 68342 107252 68348
rect 107106 68303 107162 68312
rect 107396 66978 107424 189722
rect 107488 78062 107516 190426
rect 107476 78056 107528 78062
rect 107476 77998 107528 78004
rect 107476 73772 107528 73778
rect 107476 73714 107528 73720
rect 107488 72894 107516 73714
rect 107476 72888 107528 72894
rect 107476 72830 107528 72836
rect 107580 68066 107608 199242
rect 107672 185774 107700 703582
rect 108040 703474 108068 703582
rect 108182 703520 108294 704960
rect 112046 703520 112158 704960
rect 115910 703520 116022 704960
rect 119774 703520 119886 704960
rect 123638 703520 123750 704960
rect 127502 703520 127614 704960
rect 130722 703520 130834 704960
rect 134586 703520 134698 704960
rect 138450 703520 138562 704960
rect 142314 703520 142426 704960
rect 146178 703520 146290 704960
rect 150042 703520 150154 704960
rect 153906 703520 154018 704960
rect 157770 703520 157882 704960
rect 161634 703520 161746 704960
rect 165498 703520 165610 704960
rect 169362 703520 169474 704960
rect 173226 703520 173338 704960
rect 177090 703520 177202 704960
rect 180954 703520 181066 704960
rect 184818 703520 184930 704960
rect 188038 703520 188150 704960
rect 191902 703520 192014 704960
rect 194612 703582 195652 703610
rect 108224 703474 108252 703520
rect 108040 703446 108252 703474
rect 112088 702434 112116 703520
rect 111812 702406 112116 702434
rect 111064 652792 111116 652798
rect 111064 652734 111116 652740
rect 110420 556232 110472 556238
rect 110420 556174 110472 556180
rect 109684 507884 109736 507890
rect 109684 507826 109736 507832
rect 108304 415472 108356 415478
rect 108304 415414 108356 415420
rect 108316 195906 108344 415414
rect 108396 374060 108448 374066
rect 108396 374002 108448 374008
rect 108408 197334 108436 374002
rect 108488 338156 108540 338162
rect 108488 338098 108540 338104
rect 108396 197328 108448 197334
rect 108396 197270 108448 197276
rect 108304 195900 108356 195906
rect 108304 195842 108356 195848
rect 108500 195838 108528 338098
rect 108580 309188 108632 309194
rect 108580 309130 108632 309136
rect 108488 195832 108540 195838
rect 108488 195774 108540 195780
rect 108120 192840 108172 192846
rect 108120 192782 108172 192788
rect 107660 185768 107712 185774
rect 107660 185710 107712 185716
rect 108132 136678 108160 192782
rect 108592 190534 108620 309130
rect 108672 285728 108724 285734
rect 108672 285670 108724 285676
rect 108684 195770 108712 285670
rect 108672 195764 108724 195770
rect 108672 195706 108724 195712
rect 109696 195362 109724 507826
rect 109776 491360 109828 491366
rect 109776 491302 109828 491308
rect 109684 195356 109736 195362
rect 109684 195298 109736 195304
rect 108856 195220 108908 195226
rect 108856 195162 108908 195168
rect 108672 191480 108724 191486
rect 108672 191422 108724 191428
rect 108580 190528 108632 190534
rect 108580 190470 108632 190476
rect 108580 187196 108632 187202
rect 108580 187138 108632 187144
rect 108488 185564 108540 185570
rect 108488 185506 108540 185512
rect 108396 181552 108448 181558
rect 108396 181494 108448 181500
rect 108304 148572 108356 148578
rect 108304 148514 108356 148520
rect 108210 139088 108266 139097
rect 108210 139023 108266 139032
rect 108120 136672 108172 136678
rect 108120 136614 108172 136620
rect 108224 76945 108252 139023
rect 108316 81394 108344 148514
rect 108304 81388 108356 81394
rect 108304 81330 108356 81336
rect 108316 80918 108344 81330
rect 108408 81297 108436 181494
rect 108394 81288 108450 81297
rect 108394 81223 108450 81232
rect 108304 80912 108356 80918
rect 108304 80854 108356 80860
rect 108210 76936 108266 76945
rect 108210 76871 108266 76880
rect 108500 75070 108528 185506
rect 108488 75064 108540 75070
rect 108488 75006 108540 75012
rect 108592 71738 108620 187138
rect 108684 73953 108712 191422
rect 108764 184068 108816 184074
rect 108764 184010 108816 184016
rect 108670 73944 108726 73953
rect 108670 73879 108726 73888
rect 108580 71732 108632 71738
rect 108580 71674 108632 71680
rect 107568 68060 107620 68066
rect 107568 68002 107620 68008
rect 107384 66972 107436 66978
rect 107384 66914 107436 66920
rect 108776 66774 108804 184010
rect 108868 75138 108896 195162
rect 109408 192228 109460 192234
rect 109408 192170 109460 192176
rect 109038 188592 109094 188601
rect 109038 188527 109094 188536
rect 109052 188329 109080 188527
rect 109038 188320 109094 188329
rect 109038 188255 109094 188264
rect 108948 187332 109000 187338
rect 108948 187274 109000 187280
rect 108856 75132 108908 75138
rect 108856 75074 108908 75080
rect 108960 67250 108988 187274
rect 109420 75449 109448 192170
rect 109788 191078 109816 491302
rect 109868 329860 109920 329866
rect 109868 329802 109920 329808
rect 109880 192914 109908 329802
rect 109960 260976 110012 260982
rect 109960 260918 110012 260924
rect 109972 200802 110000 260918
rect 109960 200796 110012 200802
rect 109960 200738 110012 200744
rect 110236 195492 110288 195498
rect 110236 195434 110288 195440
rect 109868 192908 109920 192914
rect 109868 192850 109920 192856
rect 109776 191072 109828 191078
rect 109776 191014 109828 191020
rect 109776 189984 109828 189990
rect 109776 189926 109828 189932
rect 109592 187740 109644 187746
rect 109592 187682 109644 187688
rect 109500 184204 109552 184210
rect 109500 184146 109552 184152
rect 109512 78849 109540 184146
rect 109498 78840 109554 78849
rect 109498 78775 109554 78784
rect 109406 75440 109462 75449
rect 109406 75375 109462 75384
rect 109604 73642 109632 187682
rect 109684 184272 109736 184278
rect 109684 184214 109736 184220
rect 109592 73636 109644 73642
rect 109592 73578 109644 73584
rect 109696 69630 109724 184214
rect 109788 74322 109816 189926
rect 110142 188320 110198 188329
rect 110142 188255 110198 188264
rect 110052 184340 110104 184346
rect 110052 184282 110104 184288
rect 109960 183932 110012 183938
rect 109960 183874 110012 183880
rect 109776 74316 109828 74322
rect 109776 74258 109828 74264
rect 109684 69624 109736 69630
rect 109684 69566 109736 69572
rect 109972 67522 110000 183874
rect 109960 67516 110012 67522
rect 109960 67458 110012 67464
rect 110064 67454 110092 184282
rect 110156 68474 110184 188255
rect 110248 72622 110276 195434
rect 110432 189038 110460 556174
rect 110512 271176 110564 271182
rect 110512 271118 110564 271124
rect 110524 270570 110552 271118
rect 110512 270564 110564 270570
rect 110512 270506 110564 270512
rect 111076 267782 111104 652734
rect 111156 369912 111208 369918
rect 111156 369854 111208 369860
rect 111064 267776 111116 267782
rect 111064 267718 111116 267724
rect 111064 262948 111116 262954
rect 111064 262890 111116 262896
rect 110420 189032 110472 189038
rect 110420 188974 110472 188980
rect 110432 187814 110460 188974
rect 110512 188760 110564 188766
rect 110512 188702 110564 188708
rect 110524 188358 110552 188702
rect 110512 188352 110564 188358
rect 110512 188294 110564 188300
rect 110420 187808 110472 187814
rect 110420 187750 110472 187756
rect 110328 184884 110380 184890
rect 110328 184826 110380 184832
rect 110236 72616 110288 72622
rect 110236 72558 110288 72564
rect 110144 68468 110196 68474
rect 110144 68410 110196 68416
rect 110052 67448 110104 67454
rect 110052 67390 110104 67396
rect 108948 67244 109000 67250
rect 108948 67186 109000 67192
rect 108764 66768 108816 66774
rect 108764 66710 108816 66716
rect 110340 52426 110368 184826
rect 110420 169040 110472 169046
rect 110420 168982 110472 168988
rect 110432 168434 110460 168982
rect 110420 168428 110472 168434
rect 110420 168370 110472 168376
rect 110696 148776 110748 148782
rect 110696 148718 110748 148724
rect 110708 71262 110736 148718
rect 110788 148232 110840 148238
rect 110788 148174 110840 148180
rect 110800 71398 110828 148174
rect 110972 144832 111024 144838
rect 110972 144774 111024 144780
rect 110880 140412 110932 140418
rect 110880 140354 110932 140360
rect 110892 72865 110920 140354
rect 110878 72856 110934 72865
rect 110878 72791 110934 72800
rect 110788 71392 110840 71398
rect 110788 71334 110840 71340
rect 110984 71330 111012 144774
rect 111076 143546 111104 262890
rect 111168 197198 111196 369854
rect 111708 270564 111760 270570
rect 111708 270506 111760 270512
rect 111340 260976 111392 260982
rect 111340 260918 111392 260924
rect 111156 197192 111208 197198
rect 111156 197134 111208 197140
rect 111156 191548 111208 191554
rect 111156 191490 111208 191496
rect 111168 190454 111196 191490
rect 111168 190426 111288 190454
rect 111260 189650 111288 190426
rect 111248 189644 111300 189650
rect 111248 189586 111300 189592
rect 111156 169040 111208 169046
rect 111156 168982 111208 168988
rect 111064 143540 111116 143546
rect 111064 143482 111116 143488
rect 111168 83473 111196 168982
rect 111154 83464 111210 83473
rect 111154 83399 111210 83408
rect 111260 79014 111288 189586
rect 111352 144362 111380 260918
rect 111524 190052 111576 190058
rect 111524 189994 111576 190000
rect 111432 188352 111484 188358
rect 111432 188294 111484 188300
rect 111340 144356 111392 144362
rect 111340 144298 111392 144304
rect 111248 79008 111300 79014
rect 111248 78950 111300 78956
rect 110972 71324 111024 71330
rect 110972 71266 111024 71272
rect 110696 71256 110748 71262
rect 110696 71198 110748 71204
rect 111444 70990 111472 188294
rect 111536 72690 111564 189994
rect 111616 187264 111668 187270
rect 111616 187206 111668 187212
rect 111524 72684 111576 72690
rect 111524 72626 111576 72632
rect 111432 70984 111484 70990
rect 111432 70926 111484 70932
rect 111628 70378 111656 187206
rect 111720 145926 111748 270506
rect 111812 200705 111840 702406
rect 115848 700528 115900 700534
rect 115848 700470 115900 700476
rect 113180 700324 113232 700330
rect 113180 700266 113232 700272
rect 111892 663808 111944 663814
rect 111892 663750 111944 663756
rect 111798 200696 111854 200705
rect 111798 200631 111854 200640
rect 111800 191276 111852 191282
rect 111800 191218 111852 191224
rect 111812 190262 111840 191218
rect 111904 191185 111932 663750
rect 112444 552084 112496 552090
rect 112444 552026 112496 552032
rect 112456 197130 112484 552026
rect 112904 263628 112956 263634
rect 112904 263570 112956 263576
rect 112536 259820 112588 259826
rect 112536 259762 112588 259768
rect 112444 197124 112496 197130
rect 112444 197066 112496 197072
rect 111984 191820 112036 191826
rect 111984 191762 112036 191768
rect 111890 191176 111946 191185
rect 111890 191111 111946 191120
rect 111800 190256 111852 190262
rect 111800 190198 111852 190204
rect 111996 190126 112024 191762
rect 111984 190120 112036 190126
rect 111984 190062 112036 190068
rect 111996 189174 112024 190062
rect 111984 189168 112036 189174
rect 111984 189110 112036 189116
rect 112444 189168 112496 189174
rect 112444 189110 112496 189116
rect 112352 186312 112404 186318
rect 112352 186254 112404 186260
rect 112168 147076 112220 147082
rect 112168 147018 112220 147024
rect 111708 145920 111760 145926
rect 111708 145862 111760 145868
rect 111708 144288 111760 144294
rect 111708 144230 111760 144236
rect 111616 70372 111668 70378
rect 111616 70314 111668 70320
rect 111720 68270 111748 144230
rect 111800 73160 111852 73166
rect 111800 73102 111852 73108
rect 111812 72350 111840 73102
rect 111800 72344 111852 72350
rect 111800 72286 111852 72292
rect 111892 68944 111944 68950
rect 111892 68886 111944 68892
rect 111708 68264 111760 68270
rect 111708 68206 111760 68212
rect 111904 68202 111932 68886
rect 111892 68196 111944 68202
rect 111892 68138 111944 68144
rect 110420 67176 110472 67182
rect 110420 67118 110472 67124
rect 110328 52420 110380 52426
rect 110328 52362 110380 52368
rect 98012 16546 98776 16574
rect 102152 16546 102640 16574
rect 106292 16546 106504 16574
rect 97816 3596 97868 3602
rect 97816 3538 97868 3544
rect 83710 354 83822 480
rect 83292 326 83822 354
rect 79846 -960 79958 326
rect 83710 -960 83822 326
rect 87574 -960 87686 480
rect 91438 -960 91550 480
rect 95302 -960 95414 480
rect 98748 354 98776 16546
rect 99166 354 99278 480
rect 98748 326 99278 354
rect 102612 354 102640 16546
rect 103030 354 103142 480
rect 102612 326 103142 354
rect 106476 354 106504 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 110432 354 110460 67118
rect 112180 65414 112208 147018
rect 112260 108316 112312 108322
rect 112260 108258 112312 108264
rect 112272 79286 112300 108258
rect 112364 80714 112392 186254
rect 112352 80708 112404 80714
rect 112352 80650 112404 80656
rect 112260 79280 112312 79286
rect 112260 79222 112312 79228
rect 112456 79150 112484 189110
rect 112548 146062 112576 259762
rect 112812 193248 112864 193254
rect 112812 193190 112864 193196
rect 112720 190256 112772 190262
rect 112720 190198 112772 190204
rect 112628 187128 112680 187134
rect 112628 187070 112680 187076
rect 112536 146056 112588 146062
rect 112536 145998 112588 146004
rect 112536 140480 112588 140486
rect 112536 140422 112588 140428
rect 112444 79144 112496 79150
rect 112444 79086 112496 79092
rect 112548 67182 112576 140422
rect 112640 72350 112668 187070
rect 112732 73030 112760 190198
rect 112824 75614 112852 193190
rect 112916 145858 112944 263570
rect 112996 262540 113048 262546
rect 112996 262482 113048 262488
rect 112904 145852 112956 145858
rect 112904 145794 112956 145800
rect 112904 145512 112956 145518
rect 112904 145454 112956 145460
rect 112812 75608 112864 75614
rect 112812 75550 112864 75556
rect 112720 73024 112772 73030
rect 112720 72966 112772 72972
rect 112628 72344 112680 72350
rect 112628 72286 112680 72292
rect 112916 69902 112944 145454
rect 113008 144226 113036 262482
rect 113192 200530 113220 700266
rect 114468 267776 114520 267782
rect 114468 267718 114520 267724
rect 114192 263900 114244 263906
rect 114192 263842 114244 263848
rect 113824 260296 113876 260302
rect 113824 260238 113876 260244
rect 113180 200524 113232 200530
rect 113180 200466 113232 200472
rect 113192 197742 113220 200466
rect 113180 197736 113232 197742
rect 113180 197678 113232 197684
rect 113088 192772 113140 192778
rect 113088 192714 113140 192720
rect 112996 144220 113048 144226
rect 112996 144162 113048 144168
rect 112904 69896 112956 69902
rect 112904 69838 112956 69844
rect 113100 68202 113128 192714
rect 113180 190528 113232 190534
rect 113180 190470 113232 190476
rect 113192 190194 113220 190470
rect 113180 190188 113232 190194
rect 113180 190130 113232 190136
rect 113732 190188 113784 190194
rect 113732 190130 113784 190136
rect 113548 153196 113600 153202
rect 113548 153138 113600 153144
rect 113560 151842 113588 153138
rect 113548 151836 113600 151842
rect 113548 151778 113600 151784
rect 113456 146124 113508 146130
rect 113456 146066 113508 146072
rect 113468 72758 113496 146066
rect 113560 80782 113588 151778
rect 113640 111852 113692 111858
rect 113640 111794 113692 111800
rect 113548 80776 113600 80782
rect 113548 80718 113600 80724
rect 113652 76294 113680 111794
rect 113744 76838 113772 190130
rect 113836 145382 113864 260238
rect 114008 259956 114060 259962
rect 114008 259898 114060 259904
rect 113916 259616 113968 259622
rect 113916 259558 113968 259564
rect 113824 145376 113876 145382
rect 113824 145318 113876 145324
rect 113928 144906 113956 259558
rect 113916 144900 113968 144906
rect 113916 144842 113968 144848
rect 114020 143177 114048 259898
rect 114100 193860 114152 193866
rect 114100 193802 114152 193808
rect 114006 143168 114062 143177
rect 114006 143103 114062 143112
rect 113824 141636 113876 141642
rect 113824 141578 113876 141584
rect 113836 79558 113864 141578
rect 114008 140616 114060 140622
rect 114008 140558 114060 140564
rect 113916 140276 113968 140282
rect 113916 140218 113968 140224
rect 113824 79552 113876 79558
rect 113824 79494 113876 79500
rect 113732 76832 113784 76838
rect 113732 76774 113784 76780
rect 113640 76288 113692 76294
rect 113640 76230 113692 76236
rect 113928 74118 113956 140218
rect 113916 74112 113968 74118
rect 113916 74054 113968 74060
rect 114020 73914 114048 140558
rect 114112 76906 114140 193802
rect 114204 145994 114232 263842
rect 114284 262404 114336 262410
rect 114284 262346 114336 262352
rect 114192 145988 114244 145994
rect 114192 145930 114244 145936
rect 114192 144900 114244 144906
rect 114192 144842 114244 144848
rect 114204 144158 114232 144842
rect 114296 144702 114324 262346
rect 114376 194472 114428 194478
rect 114376 194414 114428 194420
rect 114388 194070 114416 194414
rect 114376 194064 114428 194070
rect 114376 194006 114428 194012
rect 114284 144696 114336 144702
rect 114284 144638 114336 144644
rect 114192 144152 114244 144158
rect 114192 144094 114244 144100
rect 114284 142044 114336 142050
rect 114284 141986 114336 141992
rect 114100 76900 114152 76906
rect 114100 76842 114152 76848
rect 114008 73908 114060 73914
rect 114008 73850 114060 73856
rect 113456 72752 113508 72758
rect 113456 72694 113508 72700
rect 114296 70242 114324 141986
rect 114388 75478 114416 194006
rect 114480 144770 114508 267718
rect 115756 264036 115808 264042
rect 115756 263978 115808 263984
rect 115664 263764 115716 263770
rect 115664 263706 115716 263712
rect 115572 262472 115624 262478
rect 115572 262414 115624 262420
rect 115480 260160 115532 260166
rect 115480 260102 115532 260108
rect 115204 260024 115256 260030
rect 115204 259966 115256 259972
rect 114744 194132 114796 194138
rect 114744 194074 114796 194080
rect 114756 192302 114784 194074
rect 114928 193452 114980 193458
rect 114928 193394 114980 193400
rect 114744 192296 114796 192302
rect 114744 192238 114796 192244
rect 114836 148164 114888 148170
rect 114836 148106 114888 148112
rect 114468 144764 114520 144770
rect 114468 144706 114520 144712
rect 114744 144424 114796 144430
rect 114744 144366 114796 144372
rect 114376 75472 114428 75478
rect 114376 75414 114428 75420
rect 114756 74254 114784 144366
rect 114744 74248 114796 74254
rect 114744 74190 114796 74196
rect 114848 71670 114876 148106
rect 114940 75585 114968 193394
rect 115112 187400 115164 187406
rect 115112 187342 115164 187348
rect 115020 141704 115072 141710
rect 115020 141646 115072 141652
rect 115032 93838 115060 141646
rect 115020 93832 115072 93838
rect 115020 93774 115072 93780
rect 115032 92546 115060 93774
rect 115020 92540 115072 92546
rect 115020 92482 115072 92488
rect 115124 79626 115152 187342
rect 115216 146198 115244 259966
rect 115388 259752 115440 259758
rect 115388 259694 115440 259700
rect 115296 191276 115348 191282
rect 115296 191218 115348 191224
rect 115308 191010 115336 191218
rect 115296 191004 115348 191010
rect 115296 190946 115348 190952
rect 115204 146192 115256 146198
rect 115204 146134 115256 146140
rect 115204 143404 115256 143410
rect 115204 143346 115256 143352
rect 115216 143002 115244 143346
rect 115204 142996 115256 143002
rect 115204 142938 115256 142944
rect 115202 138952 115258 138961
rect 115202 138887 115258 138896
rect 115112 79620 115164 79626
rect 115112 79562 115164 79568
rect 115216 76566 115244 138887
rect 115308 77178 115336 190946
rect 115400 142769 115428 259694
rect 115492 143478 115520 260102
rect 115584 144634 115612 262414
rect 115572 144628 115624 144634
rect 115572 144570 115624 144576
rect 115480 143472 115532 143478
rect 115480 143414 115532 143420
rect 115676 143206 115704 263706
rect 115664 143200 115716 143206
rect 115664 143142 115716 143148
rect 115386 142760 115442 142769
rect 115386 142695 115442 142704
rect 115768 142662 115796 263978
rect 115860 190942 115888 700470
rect 115952 699854 115980 703520
rect 116032 700460 116084 700466
rect 116032 700402 116084 700408
rect 115940 699848 115992 699854
rect 115940 699790 115992 699796
rect 116044 683114 116072 700402
rect 117228 700392 117280 700398
rect 117228 700334 117280 700340
rect 115952 683086 116072 683114
rect 115952 201482 115980 683086
rect 117136 263968 117188 263974
rect 117136 263910 117188 263916
rect 116308 262608 116360 262614
rect 116308 262550 116360 262556
rect 115940 201476 115992 201482
rect 115940 201418 115992 201424
rect 115952 200394 115980 201418
rect 115940 200388 115992 200394
rect 115940 200330 115992 200336
rect 115848 190936 115900 190942
rect 115848 190878 115900 190884
rect 116216 145444 116268 145450
rect 116216 145386 116268 145392
rect 115756 142656 115808 142662
rect 115756 142598 115808 142604
rect 115572 141840 115624 141846
rect 115572 141782 115624 141788
rect 115386 140312 115442 140321
rect 115386 140247 115442 140256
rect 115296 77172 115348 77178
rect 115296 77114 115348 77120
rect 115204 76560 115256 76566
rect 115204 76502 115256 76508
rect 114926 75576 114982 75585
rect 114926 75511 114982 75520
rect 115400 73982 115428 140247
rect 115388 73976 115440 73982
rect 115388 73918 115440 73924
rect 114836 71664 114888 71670
rect 114836 71606 114888 71612
rect 114284 70236 114336 70242
rect 114284 70178 114336 70184
rect 115584 69970 115612 141782
rect 115664 141364 115716 141370
rect 115664 141306 115716 141312
rect 115572 69964 115624 69970
rect 115572 69906 115624 69912
rect 115676 69698 115704 141306
rect 115848 140548 115900 140554
rect 115848 140490 115900 140496
rect 115860 138145 115888 140490
rect 115846 138136 115902 138145
rect 115846 138071 115902 138080
rect 115846 92576 115902 92585
rect 115846 92511 115902 92520
rect 115860 81569 115888 92511
rect 115846 81560 115902 81569
rect 115846 81495 115902 81504
rect 115848 76968 115900 76974
rect 115848 76910 115900 76916
rect 115860 76566 115888 76910
rect 115848 76560 115900 76566
rect 115848 76502 115900 76508
rect 115848 69828 115900 69834
rect 115848 69770 115900 69776
rect 115860 69698 115888 69770
rect 115664 69692 115716 69698
rect 115664 69634 115716 69640
rect 115848 69692 115900 69698
rect 115848 69634 115900 69640
rect 113088 68196 113140 68202
rect 113088 68138 113140 68144
rect 112536 67176 112588 67182
rect 112536 67118 112588 67124
rect 116228 66094 116256 145386
rect 116320 143274 116348 262550
rect 116676 259888 116728 259894
rect 116676 259830 116728 259836
rect 116584 259548 116636 259554
rect 116584 259490 116636 259496
rect 116492 196444 116544 196450
rect 116492 196386 116544 196392
rect 116400 192432 116452 192438
rect 116400 192374 116452 192380
rect 116412 169046 116440 192374
rect 116504 173194 116532 196386
rect 116492 173188 116544 173194
rect 116492 173130 116544 173136
rect 116492 171828 116544 171834
rect 116492 171770 116544 171776
rect 116400 169040 116452 169046
rect 116400 168982 116452 168988
rect 116400 144492 116452 144498
rect 116400 144434 116452 144440
rect 116308 143268 116360 143274
rect 116308 143210 116360 143216
rect 116412 76265 116440 144434
rect 116398 76256 116454 76265
rect 116398 76191 116454 76200
rect 116504 66910 116532 171770
rect 116596 145625 116624 259490
rect 116688 146266 116716 259830
rect 116768 259684 116820 259690
rect 116768 259626 116820 259632
rect 116676 146260 116728 146266
rect 116676 146202 116728 146208
rect 116582 145616 116638 145625
rect 116582 145551 116638 145560
rect 116676 143268 116728 143274
rect 116676 143210 116728 143216
rect 116584 142996 116636 143002
rect 116584 142938 116636 142944
rect 116492 66904 116544 66910
rect 116492 66846 116544 66852
rect 116216 66088 116268 66094
rect 116216 66030 116268 66036
rect 112168 65408 112220 65414
rect 112168 65350 112220 65356
rect 116596 4826 116624 142938
rect 116688 142798 116716 143210
rect 116780 142934 116808 259626
rect 117044 201476 117096 201482
rect 117044 201418 117096 201424
rect 117056 198937 117084 201418
rect 117042 198928 117098 198937
rect 117042 198863 117098 198872
rect 117044 195560 117096 195566
rect 117044 195502 117096 195508
rect 116860 188760 116912 188766
rect 116860 188702 116912 188708
rect 116768 142928 116820 142934
rect 116768 142870 116820 142876
rect 116676 142792 116728 142798
rect 116676 142734 116728 142740
rect 116676 140004 116728 140010
rect 116676 139946 116728 139952
rect 116688 71466 116716 139946
rect 116768 138712 116820 138718
rect 116768 138654 116820 138660
rect 116676 71460 116728 71466
rect 116676 71402 116728 71408
rect 116780 70174 116808 138654
rect 116872 71233 116900 188702
rect 116952 155984 117004 155990
rect 116952 155926 117004 155932
rect 116964 75410 116992 155926
rect 117056 75682 117084 195502
rect 117148 142730 117176 263910
rect 117240 191554 117268 700334
rect 117964 699848 118016 699854
rect 117964 699790 118016 699796
rect 117872 259480 117924 259486
rect 117872 259422 117924 259428
rect 117320 256760 117372 256766
rect 117320 256702 117372 256708
rect 117332 200870 117360 256702
rect 117320 200864 117372 200870
rect 117320 200806 117372 200812
rect 117780 195696 117832 195702
rect 117780 195638 117832 195644
rect 117228 191548 117280 191554
rect 117228 191490 117280 191496
rect 117228 191344 117280 191350
rect 117228 191286 117280 191292
rect 117136 142724 117188 142730
rect 117136 142666 117188 142672
rect 117136 140684 117188 140690
rect 117136 140626 117188 140632
rect 117148 139505 117176 140626
rect 117134 139496 117190 139505
rect 117134 139431 117190 139440
rect 117044 75676 117096 75682
rect 117044 75618 117096 75624
rect 116952 75404 117004 75410
rect 116952 75346 117004 75352
rect 116858 71224 116914 71233
rect 116858 71159 116914 71168
rect 116768 70168 116820 70174
rect 116768 70110 116820 70116
rect 117240 66026 117268 191286
rect 117792 153202 117820 195638
rect 117780 153196 117832 153202
rect 117780 153138 117832 153144
rect 117884 145586 117912 259422
rect 117976 198966 118004 699790
rect 119816 699718 119844 703520
rect 123680 700534 123708 703520
rect 123668 700528 123720 700534
rect 123668 700470 123720 700476
rect 127544 700398 127572 703520
rect 130764 702434 130792 703520
rect 134628 702434 134656 703520
rect 138492 702434 138520 703520
rect 129936 702406 130792 702434
rect 133892 702406 134656 702434
rect 138124 702406 138520 702434
rect 127532 700392 127584 700398
rect 127532 700334 127584 700340
rect 121276 700324 121328 700330
rect 121276 700266 121328 700272
rect 119804 699712 119856 699718
rect 119804 699654 119856 699660
rect 120724 699712 120776 699718
rect 120724 699654 120776 699660
rect 120080 474768 120132 474774
rect 120080 474710 120132 474716
rect 118700 390584 118752 390590
rect 118700 390526 118752 390532
rect 118056 298172 118108 298178
rect 118056 298114 118108 298120
rect 118068 267734 118096 298114
rect 118068 267706 118188 267734
rect 118160 264994 118188 267706
rect 118148 264988 118200 264994
rect 118148 264930 118200 264936
rect 117964 198960 118016 198966
rect 117964 198902 118016 198908
rect 117964 196784 118016 196790
rect 117964 196726 118016 196732
rect 117976 181490 118004 196726
rect 118056 194132 118108 194138
rect 118056 194074 118108 194080
rect 117964 181484 118016 181490
rect 117964 181426 118016 181432
rect 117964 180260 118016 180266
rect 117964 180202 118016 180208
rect 117872 145580 117924 145586
rect 117872 145522 117924 145528
rect 117688 144560 117740 144566
rect 117688 144502 117740 144508
rect 117320 75744 117372 75750
rect 117320 75686 117372 75692
rect 117228 66020 117280 66026
rect 117228 65962 117280 65968
rect 117332 16574 117360 75686
rect 117700 71194 117728 144502
rect 117872 141500 117924 141506
rect 117872 141442 117924 141448
rect 117780 96688 117832 96694
rect 117780 96630 117832 96636
rect 117792 77042 117820 96630
rect 117780 77036 117832 77042
rect 117780 76978 117832 76984
rect 117884 75342 117912 141442
rect 117976 80646 118004 180202
rect 117964 80640 118016 80646
rect 117964 80582 118016 80588
rect 118068 79082 118096 194074
rect 118160 145722 118188 264930
rect 118516 263832 118568 263838
rect 118516 263774 118568 263780
rect 118240 262336 118292 262342
rect 118240 262278 118292 262284
rect 118148 145716 118200 145722
rect 118148 145658 118200 145664
rect 118252 142798 118280 262278
rect 118424 260840 118476 260846
rect 118424 260782 118476 260788
rect 118332 196988 118384 196994
rect 118332 196930 118384 196936
rect 118240 142792 118292 142798
rect 118240 142734 118292 142740
rect 118148 141772 118200 141778
rect 118148 141714 118200 141720
rect 118056 79076 118108 79082
rect 118056 79018 118108 79024
rect 117872 75336 117924 75342
rect 117872 75278 117924 75284
rect 118160 71641 118188 141714
rect 118240 135924 118292 135930
rect 118240 135866 118292 135872
rect 118146 71632 118202 71641
rect 118146 71567 118202 71576
rect 117688 71188 117740 71194
rect 117688 71130 117740 71136
rect 118252 70038 118280 135866
rect 118344 76770 118372 196930
rect 118436 143614 118464 260782
rect 118424 143608 118476 143614
rect 118424 143550 118476 143556
rect 118528 143138 118556 263774
rect 118712 201634 118740 390526
rect 118792 300892 118844 300898
rect 118792 300834 118844 300840
rect 118804 204354 118832 300834
rect 119988 263696 120040 263702
rect 119988 263638 120040 263644
rect 119804 262812 119856 262818
rect 119804 262754 119856 262760
rect 119620 262744 119672 262750
rect 119620 262686 119672 262692
rect 119344 252612 119396 252618
rect 119344 252554 119396 252560
rect 118804 204326 119016 204354
rect 118712 201606 118832 201634
rect 118700 201544 118752 201550
rect 118700 201486 118752 201492
rect 118712 200977 118740 201486
rect 118698 200968 118754 200977
rect 118698 200903 118754 200912
rect 118804 200462 118832 201606
rect 118988 201550 119016 204326
rect 118976 201544 119028 201550
rect 118976 201486 119028 201492
rect 119356 200598 119384 252554
rect 119436 240168 119488 240174
rect 119436 240110 119488 240116
rect 119344 200592 119396 200598
rect 119344 200534 119396 200540
rect 118792 200456 118844 200462
rect 118792 200398 118844 200404
rect 118804 200114 118832 200398
rect 119448 200114 119476 240110
rect 119528 220856 119580 220862
rect 119528 220798 119580 220804
rect 119540 200666 119568 220798
rect 119528 200660 119580 200666
rect 119528 200602 119580 200608
rect 118712 200086 118832 200114
rect 119356 200086 119476 200114
rect 118712 199617 118740 200086
rect 119356 199782 119384 200086
rect 119344 199776 119396 199782
rect 119344 199718 119396 199724
rect 118698 199608 118754 199617
rect 118698 199543 118754 199552
rect 118700 193316 118752 193322
rect 118700 193258 118752 193264
rect 118712 192370 118740 193258
rect 118700 192364 118752 192370
rect 118700 192306 118752 192312
rect 118608 191208 118660 191214
rect 118608 191150 118660 191156
rect 118516 143132 118568 143138
rect 118516 143074 118568 143080
rect 118422 138000 118478 138009
rect 118422 137935 118478 137944
rect 118332 76764 118384 76770
rect 118332 76706 118384 76712
rect 118240 70032 118292 70038
rect 118240 69974 118292 69980
rect 118436 65550 118464 137935
rect 118514 73128 118570 73137
rect 118514 73063 118570 73072
rect 118528 72894 118556 73063
rect 118516 72888 118568 72894
rect 118516 72830 118568 72836
rect 118424 65544 118476 65550
rect 118424 65486 118476 65492
rect 118620 64734 118648 191150
rect 119252 145784 119304 145790
rect 119252 145726 119304 145732
rect 119264 144974 119292 145726
rect 119068 144968 119120 144974
rect 119068 144910 119120 144916
rect 119252 144968 119304 144974
rect 119252 144910 119304 144916
rect 119080 72826 119108 144910
rect 119252 140684 119304 140690
rect 119252 140626 119304 140632
rect 119160 103556 119212 103562
rect 119160 103498 119212 103504
rect 119172 76430 119200 103498
rect 119264 80374 119292 140626
rect 119356 95198 119384 199718
rect 119436 191072 119488 191078
rect 119436 191014 119488 191020
rect 119344 95192 119396 95198
rect 119344 95134 119396 95140
rect 119344 92540 119396 92546
rect 119344 92482 119396 92488
rect 119252 80368 119304 80374
rect 119252 80310 119304 80316
rect 119356 76702 119384 92482
rect 119448 79218 119476 191014
rect 119528 189916 119580 189922
rect 119528 189858 119580 189864
rect 119436 79212 119488 79218
rect 119436 79154 119488 79160
rect 119344 76696 119396 76702
rect 119344 76638 119396 76644
rect 119160 76424 119212 76430
rect 119160 76366 119212 76372
rect 119540 74050 119568 189858
rect 119632 145654 119660 262686
rect 119712 260228 119764 260234
rect 119712 260170 119764 260176
rect 119724 191185 119752 260170
rect 119710 191176 119766 191185
rect 119710 191111 119766 191120
rect 119712 189848 119764 189854
rect 119712 189790 119764 189796
rect 119620 145648 119672 145654
rect 119620 145590 119672 145596
rect 119620 140888 119672 140894
rect 119620 140830 119672 140836
rect 119632 80442 119660 140830
rect 119620 80436 119672 80442
rect 119620 80378 119672 80384
rect 119528 74044 119580 74050
rect 119528 73986 119580 73992
rect 119540 73846 119568 73986
rect 119528 73840 119580 73846
rect 119528 73782 119580 73788
rect 119068 72820 119120 72826
rect 119068 72762 119120 72768
rect 119724 72554 119752 189790
rect 119816 142866 119844 262754
rect 119896 262676 119948 262682
rect 119896 262618 119948 262624
rect 119908 143410 119936 262618
rect 119896 143404 119948 143410
rect 119896 143346 119948 143352
rect 120000 143002 120028 263638
rect 120092 263594 120120 474710
rect 120264 289876 120316 289882
rect 120264 289818 120316 289824
rect 120092 263566 120212 263594
rect 120184 260098 120212 263566
rect 120172 260092 120224 260098
rect 120172 260034 120224 260040
rect 120080 253224 120132 253230
rect 120080 253166 120132 253172
rect 119896 142996 119948 143002
rect 119896 142938 119948 142944
rect 119988 142996 120040 143002
rect 119988 142938 120040 142944
rect 119908 142866 119936 142938
rect 120092 142866 120120 253166
rect 120184 196042 120212 260034
rect 120276 200326 120304 289818
rect 120368 259270 120612 259298
rect 120368 253230 120396 259270
rect 120356 253224 120408 253230
rect 120356 253166 120408 253172
rect 120630 218104 120686 218113
rect 120630 218039 120686 218048
rect 120540 208412 120592 208418
rect 120540 208354 120592 208360
rect 120552 200462 120580 208354
rect 120540 200456 120592 200462
rect 120540 200398 120592 200404
rect 120264 200320 120316 200326
rect 120264 200262 120316 200268
rect 120276 199170 120304 200262
rect 120264 199164 120316 199170
rect 120264 199106 120316 199112
rect 120172 196036 120224 196042
rect 120172 195978 120224 195984
rect 120356 193792 120408 193798
rect 120356 193734 120408 193740
rect 119804 142860 119856 142866
rect 119804 142802 119856 142808
rect 119896 142860 119948 142866
rect 119896 142802 119948 142808
rect 120080 142860 120132 142866
rect 120080 142802 120132 142808
rect 119816 142594 119844 142802
rect 119804 142588 119856 142594
rect 119804 142530 119856 142536
rect 119896 142112 119948 142118
rect 119896 142054 119948 142060
rect 119908 140894 119936 142054
rect 119988 141976 120040 141982
rect 119988 141918 120040 141924
rect 119896 140888 119948 140894
rect 119896 140830 119948 140836
rect 119804 139596 119856 139602
rect 119804 139538 119856 139544
rect 119816 75857 119844 139538
rect 119894 138680 119950 138689
rect 119894 138615 119950 138624
rect 119802 75848 119858 75857
rect 119802 75783 119858 75792
rect 119712 72548 119764 72554
rect 119712 72490 119764 72496
rect 119908 71602 119936 138615
rect 120000 135930 120028 141918
rect 119988 135924 120040 135930
rect 119988 135866 120040 135872
rect 120080 80912 120132 80918
rect 120080 80854 120132 80860
rect 119986 78568 120042 78577
rect 119986 78503 120042 78512
rect 120000 74186 120028 78503
rect 120092 77246 120120 80854
rect 120080 77240 120132 77246
rect 120080 77182 120132 77188
rect 120368 75002 120396 193734
rect 120644 145314 120672 218039
rect 120736 198898 120764 699654
rect 120816 503736 120868 503742
rect 120816 503678 120868 503684
rect 120724 198892 120776 198898
rect 120724 198834 120776 198840
rect 120828 198762 120856 503678
rect 121288 263594 121316 700266
rect 128360 623824 128412 623830
rect 128360 623766 128412 623772
rect 125692 608660 125744 608666
rect 125692 608602 125744 608608
rect 121460 520328 121512 520334
rect 121460 520270 121512 520276
rect 121472 267734 121500 520270
rect 124864 451308 124916 451314
rect 124864 451250 124916 451256
rect 124220 407176 124272 407182
rect 124220 407118 124272 407124
rect 122932 278044 122984 278050
rect 122932 277986 122984 277992
rect 121472 267706 121592 267734
rect 121196 263566 121316 263594
rect 121196 253934 121224 263566
rect 121564 262886 121592 267706
rect 122944 263594 122972 277986
rect 124232 267734 124260 407118
rect 124232 267706 124352 267734
rect 124324 263594 124352 267706
rect 124876 264042 124904 451250
rect 125704 267734 125732 608602
rect 126980 313336 127032 313342
rect 126980 313278 127032 313284
rect 125704 267706 126008 267734
rect 124864 264036 124916 264042
rect 124864 263978 124916 263984
rect 125232 264036 125284 264042
rect 125232 263978 125284 263984
rect 122944 263566 123248 263594
rect 124324 263566 124444 263594
rect 121552 262880 121604 262886
rect 121552 262822 121604 262828
rect 121564 262313 121592 262822
rect 122562 262712 122618 262721
rect 122562 262647 122618 262656
rect 121550 262304 121606 262313
rect 121550 262239 121606 262248
rect 121368 260092 121420 260098
rect 121368 260034 121420 260040
rect 121380 259978 121408 260034
rect 122576 260001 122604 262647
rect 122840 260840 122892 260846
rect 122840 260782 122892 260788
rect 122562 259992 122618 260001
rect 121380 259950 121440 259978
rect 122268 259950 122562 259978
rect 122852 259978 122880 260782
rect 122852 259950 123096 259978
rect 123220 259962 123248 263566
rect 124416 260302 124444 263566
rect 124404 260296 124456 260302
rect 124404 260238 124456 260244
rect 124416 259978 124444 260238
rect 125244 259978 125272 263978
rect 125980 263594 126008 267706
rect 126992 263974 127020 313278
rect 128372 267734 128400 623766
rect 128372 267706 128492 267734
rect 126980 263968 127032 263974
rect 126980 263910 127032 263916
rect 127716 263968 127768 263974
rect 127716 263910 127768 263916
rect 125980 263566 126100 263594
rect 126072 260030 126100 263566
rect 126980 262948 127032 262954
rect 126980 262890 127032 262896
rect 126060 260024 126112 260030
rect 123588 259962 123924 259978
rect 123208 259956 123260 259962
rect 122562 259927 122618 259936
rect 122576 259867 122604 259927
rect 123208 259898 123260 259904
rect 123576 259956 123924 259962
rect 123628 259950 123924 259956
rect 124416 259950 124752 259978
rect 125244 259950 125580 259978
rect 126992 259978 127020 262890
rect 127728 259978 127756 263910
rect 128464 259978 128492 267706
rect 129936 260846 129964 702406
rect 131120 467900 131172 467906
rect 131120 467842 131172 467848
rect 130016 263084 130068 263090
rect 130016 263026 130068 263032
rect 129740 260840 129792 260846
rect 129740 260782 129792 260788
rect 129924 260840 129976 260846
rect 129924 260782 129976 260788
rect 129752 260166 129780 260782
rect 129740 260160 129792 260166
rect 129740 260102 129792 260108
rect 126112 259972 126408 259978
rect 126060 259966 126408 259972
rect 126072 259950 126408 259966
rect 126992 259950 127236 259978
rect 127728 259950 128064 259978
rect 128464 259950 128892 259978
rect 123576 259898 123628 259904
rect 128464 259894 128492 259950
rect 128452 259888 128504 259894
rect 128452 259830 128504 259836
rect 129370 259720 129426 259729
rect 130028 259706 130056 263026
rect 130200 262336 130252 262342
rect 130200 262278 130252 262284
rect 130212 259978 130240 262278
rect 130212 259950 130548 259978
rect 131132 259842 131160 467842
rect 132592 269816 132644 269822
rect 132592 269758 132644 269764
rect 132604 263906 132632 269758
rect 133892 265810 133920 702406
rect 133972 270564 134024 270570
rect 133972 270506 134024 270512
rect 133984 267734 134012 270506
rect 133984 267706 134288 267734
rect 133880 265804 133932 265810
rect 133880 265746 133932 265752
rect 132592 263900 132644 263906
rect 132592 263842 132644 263848
rect 133512 263900 133564 263906
rect 133512 263842 133564 263848
rect 132132 263560 132184 263566
rect 132132 263502 132184 263508
rect 131132 259826 131376 259842
rect 131120 259820 131376 259826
rect 131172 259814 131376 259820
rect 131120 259762 131172 259768
rect 132144 259706 132172 263502
rect 132684 260840 132736 260846
rect 132684 260782 132736 260788
rect 132696 259978 132724 260782
rect 133524 259978 133552 263842
rect 134260 259978 134288 267706
rect 136548 265736 136600 265742
rect 136548 265678 136600 265684
rect 136560 263809 136588 265678
rect 135442 263800 135498 263809
rect 135442 263735 135498 263744
rect 136546 263800 136602 263809
rect 136546 263735 136602 263744
rect 134890 262848 134946 262857
rect 134890 262783 134946 262792
rect 134904 262274 134932 262783
rect 134892 262268 134944 262274
rect 134892 262210 134944 262216
rect 132696 259950 133032 259978
rect 133524 259950 133860 259978
rect 134260 259950 134688 259978
rect 135456 259842 135484 263735
rect 137652 262676 137704 262682
rect 137652 262618 137704 262624
rect 136824 262540 136876 262546
rect 136824 262482 136876 262488
rect 135996 262268 136048 262274
rect 135996 262210 136048 262216
rect 136008 259978 136036 262210
rect 136836 259978 136864 262482
rect 137664 259978 137692 262618
rect 138124 260137 138152 702406
rect 142356 683114 142384 703520
rect 146220 697610 146248 703520
rect 150084 702434 150112 703520
rect 153948 702434 153976 703520
rect 149072 702406 150112 702434
rect 153212 702406 153976 702434
rect 144920 697604 144972 697610
rect 144920 697546 144972 697552
rect 146208 697604 146260 697610
rect 146208 697546 146260 697552
rect 142172 683086 142384 683114
rect 139492 267776 139544 267782
rect 139492 267718 139544 267724
rect 138480 262880 138532 262886
rect 138480 262822 138532 262828
rect 138110 260128 138166 260137
rect 138110 260063 138166 260072
rect 138492 259978 138520 262822
rect 139504 259978 139532 267718
rect 140780 262948 140832 262954
rect 140780 262890 140832 262896
rect 140136 262608 140188 262614
rect 140136 262550 140188 262556
rect 140148 259978 140176 262550
rect 140792 262410 140820 262890
rect 141792 262472 141844 262478
rect 141792 262414 141844 262420
rect 140780 262404 140832 262410
rect 140780 262346 140832 262352
rect 140792 260148 140820 262346
rect 140792 260120 140912 260148
rect 140884 259978 140912 260120
rect 141804 259978 141832 262414
rect 142172 260166 142200 683086
rect 142804 271176 142856 271182
rect 142804 271118 142856 271124
rect 142816 267734 142844 271118
rect 142632 267706 142844 267734
rect 142632 263770 142660 267706
rect 144828 267096 144880 267102
rect 144828 267038 144880 267044
rect 142620 263764 142672 263770
rect 142620 263706 142672 263712
rect 142160 260160 142212 260166
rect 142160 260102 142212 260108
rect 142632 259978 142660 263706
rect 144840 263634 144868 267038
rect 143724 263628 143776 263634
rect 143724 263570 143776 263576
rect 144828 263628 144880 263634
rect 144828 263570 144880 263576
rect 136008 259950 136344 259978
rect 136836 259950 137172 259978
rect 137664 259950 138000 259978
rect 138492 259950 138828 259978
rect 139504 259950 139656 259978
rect 140148 259950 140484 259978
rect 140884 259950 141312 259978
rect 141804 259950 142140 259978
rect 142632 259950 142968 259978
rect 143736 259842 143764 263570
rect 144828 260976 144880 260982
rect 144828 260918 144880 260924
rect 144840 259978 144868 260918
rect 144932 260234 144960 697546
rect 147680 273964 147732 273970
rect 147680 273906 147732 273912
rect 145012 268388 145064 268394
rect 145012 268330 145064 268336
rect 145024 260234 145052 268330
rect 146208 264444 146260 264450
rect 146208 264386 146260 264392
rect 146220 263838 146248 264386
rect 145380 263832 145432 263838
rect 145380 263774 145432 263780
rect 146208 263832 146260 263838
rect 146208 263774 146260 263780
rect 144920 260228 144972 260234
rect 144920 260170 144972 260176
rect 145012 260228 145064 260234
rect 145012 260170 145064 260176
rect 144624 259950 144868 259978
rect 135456 259814 135516 259842
rect 143736 259814 143796 259842
rect 145024 259758 145052 260170
rect 145392 259842 145420 263774
rect 147692 260234 147720 273906
rect 148048 265668 148100 265674
rect 148048 265610 148100 265616
rect 148060 263945 148088 265610
rect 148046 263936 148102 263945
rect 148046 263871 148102 263880
rect 146254 260228 146306 260234
rect 146254 260170 146306 260176
rect 147680 260228 147732 260234
rect 147680 260170 147732 260176
rect 146266 259964 146294 260170
rect 145392 259814 145452 259842
rect 145012 259752 145064 259758
rect 129426 259678 130056 259706
rect 131868 259678 132204 259706
rect 145012 259694 145064 259700
rect 147692 259690 147720 260170
rect 148060 259842 148088 263871
rect 149072 260234 149100 702406
rect 149152 271244 149204 271250
rect 149152 271186 149204 271192
rect 148738 260228 148790 260234
rect 148738 260170 148790 260176
rect 149060 260228 149112 260234
rect 149060 260170 149112 260176
rect 148750 259964 148778 260170
rect 149164 259978 149192 271186
rect 153212 265878 153240 702406
rect 157812 700330 157840 703520
rect 157800 700324 157852 700330
rect 157800 700266 157852 700272
rect 161676 683114 161704 703520
rect 165540 700398 165568 703520
rect 169404 700466 169432 703520
rect 177132 700534 177160 703520
rect 177120 700528 177172 700534
rect 177120 700470 177172 700476
rect 169392 700460 169444 700466
rect 169392 700402 169444 700408
rect 165528 700392 165580 700398
rect 165528 700334 165580 700340
rect 180996 700126 181024 703520
rect 184860 700670 184888 703520
rect 184848 700664 184900 700670
rect 184848 700606 184900 700612
rect 188080 700602 188108 703520
rect 188068 700596 188120 700602
rect 188068 700538 188120 700544
rect 191840 700460 191892 700466
rect 191840 700402 191892 700408
rect 194508 700460 194560 700466
rect 194508 700402 194560 700408
rect 189724 700324 189776 700330
rect 189724 700266 189776 700272
rect 180984 700120 181036 700126
rect 180984 700062 181036 700068
rect 189448 700120 189500 700126
rect 189448 700062 189500 700068
rect 181444 684548 181496 684554
rect 181444 684490 181496 684496
rect 161492 683086 161704 683114
rect 155960 271924 156012 271930
rect 155960 271866 156012 271872
rect 153200 265872 153252 265878
rect 153200 265814 153252 265820
rect 151912 264988 151964 264994
rect 151912 264930 151964 264936
rect 154488 264988 154540 264994
rect 154488 264930 154540 264936
rect 149244 264240 149296 264246
rect 149244 264182 149296 264188
rect 150348 264240 150400 264246
rect 150348 264182 150400 264188
rect 149256 263702 149284 264182
rect 149244 263696 149296 263702
rect 149244 263638 149296 263644
rect 150360 259978 150388 264182
rect 151924 259978 151952 264930
rect 152556 262812 152608 262818
rect 152556 262754 152608 262760
rect 152568 259978 152596 262754
rect 153384 262744 153436 262750
rect 153384 262686 153436 262692
rect 153396 259978 153424 262686
rect 154500 259978 154528 264930
rect 155684 262812 155736 262818
rect 155684 262754 155736 262760
rect 155696 259978 155724 262754
rect 147936 259814 148088 259842
rect 149164 259950 149592 259978
rect 150360 259950 150420 259978
rect 151924 259950 152076 259978
rect 152568 259950 152904 259978
rect 153396 259950 153732 259978
rect 154500 259950 154560 259978
rect 155388 259950 155724 259978
rect 155972 259978 156000 271866
rect 160100 268456 160152 268462
rect 160100 268398 160152 268404
rect 158720 264376 158772 264382
rect 158720 264318 158772 264324
rect 158352 264308 158404 264314
rect 158352 264250 158404 264256
rect 157248 263152 157300 263158
rect 157248 263094 157300 263100
rect 157260 259978 157288 263094
rect 158168 262404 158220 262410
rect 158168 262346 158220 262352
rect 158180 259978 158208 262346
rect 158364 260302 158392 264250
rect 158732 263634 158760 264318
rect 158720 263628 158772 263634
rect 158720 263570 158772 263576
rect 159456 263628 159508 263634
rect 159456 263570 159508 263576
rect 158352 260296 158404 260302
rect 158352 260238 158404 260244
rect 155972 259950 156216 259978
rect 157044 259950 157288 259978
rect 157872 259950 158208 259978
rect 158364 259978 158392 260238
rect 159468 259978 159496 263570
rect 160112 260098 160140 268398
rect 161492 265946 161520 683086
rect 179420 398880 179472 398886
rect 179420 398822 179472 398828
rect 178040 354748 178092 354754
rect 178040 354690 178092 354696
rect 170404 294024 170456 294030
rect 170404 293966 170456 293972
rect 169760 276072 169812 276078
rect 169760 276014 169812 276020
rect 169772 267734 169800 276014
rect 169772 267706 170352 267734
rect 167460 267028 167512 267034
rect 167460 266970 167512 266976
rect 163964 266416 164016 266422
rect 163964 266358 164016 266364
rect 161480 265940 161532 265946
rect 161480 265882 161532 265888
rect 161940 263424 161992 263430
rect 161940 263366 161992 263372
rect 160652 262472 160704 262478
rect 160652 262414 160704 262420
rect 160100 260092 160152 260098
rect 160100 260034 160152 260040
rect 160664 259978 160692 262414
rect 161204 260364 161256 260370
rect 161204 260306 161256 260312
rect 161216 260250 161244 260306
rect 161170 260222 161244 260250
rect 161170 260098 161198 260222
rect 161158 260092 161210 260098
rect 161158 260034 161210 260040
rect 158364 259950 158700 259978
rect 159468 259950 159528 259978
rect 160356 259950 160692 259978
rect 161170 259964 161198 260034
rect 147680 259684 147732 259690
rect 129370 259655 129426 259664
rect 131868 259593 131896 259678
rect 147680 259626 147732 259632
rect 146760 259616 146812 259622
rect 131854 259584 131910 259593
rect 146812 259564 147108 259570
rect 146760 259558 147108 259564
rect 146772 259542 147108 259558
rect 149164 259554 149192 259950
rect 161952 259570 161980 263366
rect 162768 261044 162820 261050
rect 162768 260986 162820 260992
rect 162780 259978 162808 260986
rect 163976 259978 164004 266358
rect 166724 263764 166776 263770
rect 166724 263706 166776 263712
rect 166736 263498 166764 263706
rect 166724 263492 166776 263498
rect 166724 263434 166776 263440
rect 164792 262880 164844 262886
rect 164792 262822 164844 262828
rect 164804 259978 164832 262822
rect 165528 262540 165580 262546
rect 165528 262482 165580 262488
rect 165540 259978 165568 262482
rect 162780 259950 162840 259978
rect 163668 259950 164004 259978
rect 164496 259950 164832 259978
rect 165324 259950 165568 259978
rect 166736 259978 166764 263434
rect 167472 259978 167500 266970
rect 169760 266484 169812 266490
rect 169760 266426 169812 266432
rect 168930 263664 168986 263673
rect 169772 263650 169800 266426
rect 168930 263599 168986 263608
rect 169680 263622 169800 263650
rect 168944 259978 168972 263599
rect 169680 259978 169708 263622
rect 170324 262834 170352 267706
rect 170416 267102 170444 293966
rect 170404 267096 170456 267102
rect 170404 267038 170456 267044
rect 171600 263356 171652 263362
rect 171600 263298 171652 263304
rect 170324 262806 170720 262834
rect 170588 262744 170640 262750
rect 170588 262686 170640 262692
rect 170600 259978 170628 262686
rect 166736 259950 166980 259978
rect 167472 259950 167960 259978
rect 168636 259950 168972 259978
rect 169464 259950 169708 259978
rect 170292 259950 170628 259978
rect 170692 259978 170720 262806
rect 170692 259950 171120 259978
rect 167932 259826 167960 259950
rect 167920 259820 167972 259826
rect 167920 259762 167972 259768
rect 171612 259706 171640 263298
rect 174728 262676 174780 262682
rect 174728 262618 174780 262624
rect 173808 262608 173860 262614
rect 173808 262550 173860 262556
rect 173072 262268 173124 262274
rect 173072 262210 173124 262216
rect 173084 259978 173112 262210
rect 173820 259978 173848 262550
rect 174740 259978 174768 262618
rect 177948 262336 178000 262342
rect 177948 262278 178000 262284
rect 176660 260908 176712 260914
rect 176660 260850 176712 260856
rect 172776 259950 173112 259978
rect 173604 259950 173848 259978
rect 174432 259950 174768 259978
rect 176672 259978 176700 260850
rect 177960 259978 177988 262278
rect 178052 260098 178080 354690
rect 179432 267734 179460 398822
rect 179432 267706 179828 267734
rect 179418 262848 179474 262857
rect 179418 262783 179474 262792
rect 179432 262342 179460 262783
rect 179420 262336 179472 262342
rect 179420 262278 179472 262284
rect 178040 260092 178092 260098
rect 178040 260034 178092 260040
rect 179374 260092 179426 260098
rect 179374 260034 179426 260040
rect 179386 259978 179414 260034
rect 179800 259978 179828 267706
rect 181456 262449 181484 684490
rect 182180 483064 182232 483070
rect 182180 483006 182232 483012
rect 181442 262440 181498 262449
rect 181442 262375 181498 262384
rect 181352 262336 181404 262342
rect 181352 262278 181404 262284
rect 180340 260024 180392 260030
rect 176672 259950 176916 259978
rect 177744 259950 177988 259978
rect 178572 259962 178908 259978
rect 179386 259964 179552 259978
rect 178572 259956 178920 259962
rect 178572 259950 178868 259956
rect 179400 259950 179552 259964
rect 179800 259972 180340 259978
rect 181364 259978 181392 262278
rect 179800 259966 180392 259972
rect 179800 259950 180380 259966
rect 181056 259950 181392 259978
rect 181456 259978 181484 262375
rect 182192 260001 182220 483006
rect 184940 375420 184992 375426
rect 184940 375362 184992 375368
rect 183652 269136 183704 269142
rect 183652 269078 183704 269084
rect 183664 267734 183692 269078
rect 183664 267706 183968 267734
rect 183006 262984 183062 262993
rect 183006 262919 183062 262928
rect 182178 259992 182234 260001
rect 181456 259950 181884 259978
rect 178868 259898 178920 259904
rect 179524 259894 179552 259950
rect 183020 259978 183048 262919
rect 182712 259950 183048 259978
rect 183374 259992 183430 260001
rect 182178 259927 182234 259936
rect 183940 259978 183968 267706
rect 184664 260024 184716 260030
rect 183430 259950 183540 259978
rect 183940 259972 184664 259978
rect 184952 260001 184980 375362
rect 189080 266008 189132 266014
rect 189080 265950 189132 265956
rect 189092 264994 189120 265950
rect 189080 264988 189132 264994
rect 189080 264930 189132 264936
rect 185490 262576 185546 262585
rect 185490 262511 185546 262520
rect 183940 259966 184716 259972
rect 184938 259992 184994 260001
rect 183940 259950 184704 259966
rect 183374 259927 183430 259936
rect 185504 259978 185532 262511
rect 185196 259950 185532 259978
rect 185858 259992 185914 260001
rect 184938 259927 184994 259936
rect 185914 259950 186024 259978
rect 185858 259927 185914 259936
rect 179512 259888 179564 259894
rect 179512 259830 179564 259836
rect 172244 259752 172296 259758
rect 166152 259690 166488 259706
rect 171612 259700 172244 259706
rect 171612 259694 172296 259700
rect 166152 259684 166500 259690
rect 166152 259678 166448 259684
rect 171612 259678 172284 259694
rect 166448 259626 166500 259632
rect 162308 259616 162360 259622
rect 149152 259548 149204 259554
rect 131854 259519 131910 259528
rect 149152 259490 149204 259496
rect 150912 259542 151248 259570
rect 161952 259564 162308 259570
rect 183388 259593 183416 259927
rect 183374 259584 183430 259593
rect 161952 259558 162360 259564
rect 161952 259542 162348 259558
rect 175260 259554 175412 259570
rect 175260 259548 175424 259554
rect 175260 259542 175372 259548
rect 150912 259486 150940 259542
rect 176088 259542 176424 259570
rect 175372 259490 175424 259496
rect 176396 259486 176424 259542
rect 183374 259519 183430 259528
rect 150900 259480 150952 259486
rect 150900 259422 150952 259428
rect 176384 259480 176436 259486
rect 176384 259422 176436 259428
rect 186962 259312 187018 259321
rect 186852 259270 186962 259298
rect 186962 259247 187018 259256
rect 121196 253906 121316 253934
rect 120908 229152 120960 229158
rect 120908 229094 120960 229100
rect 120920 198830 120948 229094
rect 121184 200796 121236 200802
rect 121184 200738 121236 200744
rect 121196 200530 121224 200738
rect 121184 200524 121236 200530
rect 121184 200466 121236 200472
rect 121000 200456 121052 200462
rect 121000 200398 121052 200404
rect 121012 199850 121040 200398
rect 121000 199844 121052 199850
rect 121000 199786 121052 199792
rect 121288 199374 121316 253906
rect 125554 200728 125606 200734
rect 122838 200696 122894 200705
rect 125692 200728 125744 200734
rect 125606 200676 125640 200682
rect 125554 200670 125640 200676
rect 125692 200670 125744 200676
rect 129002 200696 129058 200705
rect 125566 200654 125640 200670
rect 122838 200631 122894 200640
rect 121276 199368 121328 199374
rect 121276 199310 121328 199316
rect 120908 198824 120960 198830
rect 120908 198766 120960 198772
rect 120816 198756 120868 198762
rect 120816 198698 120868 198704
rect 120724 198688 120776 198694
rect 120724 198630 120776 198636
rect 120736 180985 120764 198630
rect 121184 198620 121236 198626
rect 121184 198562 121236 198568
rect 121092 184476 121144 184482
rect 121092 184418 121144 184424
rect 120722 180976 120778 180985
rect 120722 180911 120778 180920
rect 120736 180538 120764 180911
rect 120724 180532 120776 180538
rect 120724 180474 120776 180480
rect 121000 180328 121052 180334
rect 121000 180270 121052 180276
rect 120908 176044 120960 176050
rect 120908 175986 120960 175992
rect 120816 148300 120868 148306
rect 120816 148242 120868 148248
rect 120632 145308 120684 145314
rect 120632 145250 120684 145256
rect 120448 143200 120500 143206
rect 120500 143148 120672 143154
rect 120448 143142 120672 143148
rect 120460 143126 120672 143142
rect 120644 143070 120672 143126
rect 120632 143064 120684 143070
rect 120632 143006 120684 143012
rect 120630 139088 120686 139097
rect 120630 139023 120686 139032
rect 120540 95192 120592 95198
rect 120540 95134 120592 95140
rect 120356 74996 120408 75002
rect 120356 74938 120408 74944
rect 120552 74390 120580 95134
rect 120540 74384 120592 74390
rect 120540 74326 120592 74332
rect 119988 74180 120040 74186
rect 119988 74122 120040 74128
rect 119896 71596 119948 71602
rect 119896 71538 119948 71544
rect 120644 70106 120672 139023
rect 120722 138544 120778 138553
rect 120722 138479 120778 138488
rect 120736 70310 120764 138479
rect 120724 70304 120776 70310
rect 120724 70246 120776 70252
rect 120632 70100 120684 70106
rect 120632 70042 120684 70048
rect 120828 66230 120856 148242
rect 120920 80918 120948 175986
rect 120908 80912 120960 80918
rect 120908 80854 120960 80860
rect 121012 78674 121040 180270
rect 121000 78668 121052 78674
rect 121000 78610 121052 78616
rect 121104 75750 121132 184418
rect 121196 79422 121224 198562
rect 121288 198558 121316 199310
rect 121276 198552 121328 198558
rect 121276 198494 121328 198500
rect 122196 197940 122248 197946
rect 122196 197882 122248 197888
rect 121276 196580 121328 196586
rect 121276 196522 121328 196528
rect 121184 79416 121236 79422
rect 121184 79358 121236 79364
rect 121288 78198 121316 196522
rect 121460 196036 121512 196042
rect 121460 195978 121512 195984
rect 121366 194576 121422 194585
rect 121366 194511 121422 194520
rect 121380 194138 121408 194511
rect 121368 194132 121420 194138
rect 121368 194074 121420 194080
rect 121368 145308 121420 145314
rect 121368 145250 121420 145256
rect 121380 143342 121408 145250
rect 121472 143546 121500 195978
rect 122104 195628 122156 195634
rect 122104 195570 122156 195576
rect 122012 193724 122064 193730
rect 122012 193666 122064 193672
rect 121552 186176 121604 186182
rect 121552 186118 121604 186124
rect 121564 185502 121592 186118
rect 121552 185496 121604 185502
rect 121552 185438 121604 185444
rect 121920 185496 121972 185502
rect 121920 185438 121972 185444
rect 121828 144900 121880 144906
rect 121828 144842 121880 144848
rect 121552 143676 121604 143682
rect 121552 143618 121604 143624
rect 121460 143540 121512 143546
rect 121460 143482 121512 143488
rect 121564 143410 121592 143618
rect 121552 143404 121604 143410
rect 121552 143346 121604 143352
rect 121368 143336 121420 143342
rect 121368 143278 121420 143284
rect 121368 142860 121420 142866
rect 121368 142802 121420 142808
rect 121380 139890 121408 142802
rect 121380 139862 121440 139890
rect 121734 122768 121790 122777
rect 121734 122703 121790 122712
rect 121748 113257 121776 122703
rect 121734 113248 121790 113257
rect 121734 113183 121790 113192
rect 121734 113112 121790 113121
rect 121734 113047 121790 113056
rect 121748 103601 121776 113047
rect 121734 103592 121790 103601
rect 121734 103527 121790 103536
rect 121734 103456 121790 103465
rect 121734 103391 121790 103400
rect 121748 93945 121776 103391
rect 121734 93936 121790 93945
rect 121734 93871 121790 93880
rect 121734 93800 121790 93809
rect 121734 93735 121790 93744
rect 121276 78192 121328 78198
rect 121276 78134 121328 78140
rect 121092 75744 121144 75750
rect 121092 75686 121144 75692
rect 121748 68950 121776 93735
rect 121736 68944 121788 68950
rect 121736 68886 121788 68892
rect 120816 66224 120868 66230
rect 120816 66166 120868 66172
rect 121840 65278 121868 144842
rect 121932 78946 121960 185438
rect 121920 78940 121972 78946
rect 121920 78882 121972 78888
rect 122024 77722 122052 193666
rect 122012 77716 122064 77722
rect 122012 77658 122064 77664
rect 121828 65272 121880 65278
rect 121828 65214 121880 65220
rect 118608 64728 118660 64734
rect 118608 64670 118660 64676
rect 122116 64394 122144 195570
rect 122208 176730 122236 197882
rect 122852 197441 122880 200631
rect 124404 200524 124456 200530
rect 124404 200466 124456 200472
rect 123206 200424 123262 200433
rect 123206 200359 123262 200368
rect 123220 200326 123248 200359
rect 123208 200320 123260 200326
rect 123208 200262 123260 200268
rect 122838 197432 122894 197441
rect 122838 197367 122894 197376
rect 122838 195936 122894 195945
rect 122838 195871 122894 195880
rect 122196 176724 122248 176730
rect 122196 176666 122248 176672
rect 122196 143540 122248 143546
rect 122196 143482 122248 143488
rect 122288 143540 122340 143546
rect 122288 143482 122340 143488
rect 122208 139890 122236 143482
rect 122300 143274 122328 143482
rect 122288 143268 122340 143274
rect 122288 143210 122340 143216
rect 122288 142860 122340 142866
rect 122288 142802 122340 142808
rect 122300 142594 122328 142802
rect 122288 142588 122340 142594
rect 122288 142530 122340 142536
rect 122852 139890 122880 195871
rect 122932 188896 122984 188902
rect 122932 188838 122984 188844
rect 122944 145450 122972 188838
rect 122932 145444 122984 145450
rect 122932 145386 122984 145392
rect 123220 140690 123248 200262
rect 124312 198892 124364 198898
rect 124312 198834 124364 198840
rect 124126 198248 124182 198257
rect 124126 198183 124182 198192
rect 124140 197441 124168 198183
rect 124126 197432 124182 197441
rect 124126 197367 124182 197376
rect 123482 193896 123538 193905
rect 123482 193831 123538 193840
rect 123496 179489 123524 193831
rect 124034 192536 124090 192545
rect 124034 192471 124090 192480
rect 123760 188896 123812 188902
rect 123760 188838 123812 188844
rect 123772 188290 123800 188838
rect 123760 188284 123812 188290
rect 123760 188226 123812 188232
rect 124048 180674 124076 192471
rect 124036 180668 124088 180674
rect 124036 180610 124088 180616
rect 124048 179602 124076 180610
rect 123956 179574 124076 179602
rect 123482 179480 123538 179489
rect 123482 179415 123538 179424
rect 123956 171134 123984 179574
rect 124034 179480 124090 179489
rect 124034 179415 124090 179424
rect 124048 179110 124076 179415
rect 124036 179104 124088 179110
rect 124036 179046 124088 179052
rect 123956 171106 124076 171134
rect 123668 143608 123720 143614
rect 123668 143550 123720 143556
rect 123208 140684 123260 140690
rect 123208 140626 123260 140632
rect 123484 140208 123536 140214
rect 123484 140150 123536 140156
rect 123496 140010 123524 140150
rect 123484 140004 123536 140010
rect 123484 139946 123536 139952
rect 123680 139890 123708 143550
rect 122208 139862 122268 139890
rect 122852 139862 123096 139890
rect 123680 139862 123924 139890
rect 124048 139369 124076 171106
rect 124140 139505 124168 197367
rect 124220 192500 124272 192506
rect 124220 192442 124272 192448
rect 124232 145518 124260 192442
rect 124220 145512 124272 145518
rect 124220 145454 124272 145460
rect 124324 139913 124352 198834
rect 124416 196722 124444 200466
rect 125612 199073 125640 200654
rect 125704 199102 125732 200670
rect 129002 200631 129058 200640
rect 177948 200660 178000 200666
rect 127162 199880 127218 199889
rect 127162 199815 127218 199824
rect 127900 199844 127952 199850
rect 126150 199744 126206 199753
rect 126150 199679 126206 199688
rect 125692 199096 125744 199102
rect 125598 199064 125654 199073
rect 125692 199038 125744 199044
rect 125598 198999 125654 199008
rect 125508 198892 125560 198898
rect 125508 198834 125560 198840
rect 125520 198762 125548 198834
rect 124772 198756 124824 198762
rect 124772 198698 124824 198704
rect 125508 198756 125560 198762
rect 125508 198698 125560 198704
rect 124784 197713 124812 198698
rect 126164 198218 126192 199679
rect 126520 198688 126572 198694
rect 126520 198630 126572 198636
rect 126532 198422 126560 198630
rect 126520 198416 126572 198422
rect 126520 198358 126572 198364
rect 126152 198212 126204 198218
rect 126152 198154 126204 198160
rect 126886 198112 126942 198121
rect 126886 198047 126942 198056
rect 124770 197704 124826 197713
rect 124770 197639 124826 197648
rect 124404 196716 124456 196722
rect 124404 196658 124456 196664
rect 124784 190454 124812 197639
rect 125506 197568 125562 197577
rect 125506 197503 125562 197512
rect 125414 197160 125470 197169
rect 125414 197095 125470 197104
rect 125428 196586 125456 197095
rect 125416 196580 125468 196586
rect 125416 196522 125468 196528
rect 124956 193248 125008 193254
rect 124956 193190 125008 193196
rect 124784 190426 124904 190454
rect 124770 179616 124826 179625
rect 124770 179551 124826 179560
rect 124784 179178 124812 179551
rect 124772 179172 124824 179178
rect 124772 179114 124824 179120
rect 124402 143168 124458 143177
rect 124402 143103 124458 143112
rect 124310 139904 124366 139913
rect 124416 139890 124444 143103
rect 124876 140622 124904 190426
rect 124864 140616 124916 140622
rect 124864 140558 124916 140564
rect 124416 139862 124752 139890
rect 124310 139839 124366 139848
rect 124968 139602 124996 193190
rect 125520 192506 125548 197503
rect 125508 192500 125560 192506
rect 125508 192442 125560 192448
rect 126796 188828 126848 188834
rect 126796 188770 126848 188776
rect 126808 187474 126836 188770
rect 126244 187468 126296 187474
rect 126244 187410 126296 187416
rect 126796 187468 126848 187474
rect 126796 187410 126848 187416
rect 125692 182844 125744 182850
rect 125692 182786 125744 182792
rect 125704 151814 125732 182786
rect 126256 151814 126284 187410
rect 126900 181490 126928 198047
rect 127176 198014 127204 199815
rect 127900 199786 127952 199792
rect 127714 198520 127770 198529
rect 127714 198455 127770 198464
rect 127164 198008 127216 198014
rect 127164 197950 127216 197956
rect 126978 194304 127034 194313
rect 126978 194239 127034 194248
rect 126992 194002 127020 194239
rect 126980 193996 127032 194002
rect 126980 193938 127032 193944
rect 127624 192500 127676 192506
rect 127624 192442 127676 192448
rect 126888 181484 126940 181490
rect 126888 181426 126940 181432
rect 126900 180794 126928 181426
rect 126900 180766 127020 180794
rect 125704 151786 125916 151814
rect 125232 145376 125284 145382
rect 125232 145318 125284 145324
rect 125244 139890 125272 145318
rect 125244 139862 125580 139890
rect 125888 139641 125916 151786
rect 125980 151786 126284 151814
rect 125874 139632 125930 139641
rect 124956 139596 125008 139602
rect 125874 139567 125930 139576
rect 124956 139538 125008 139544
rect 124126 139496 124182 139505
rect 124126 139431 124182 139440
rect 125980 139369 126008 151786
rect 126992 148617 127020 180766
rect 127636 155922 127664 192442
rect 127728 179761 127756 198455
rect 127808 197804 127860 197810
rect 127808 197746 127860 197752
rect 127820 180878 127848 197746
rect 127912 192545 127940 199786
rect 128452 199572 128504 199578
rect 128452 199514 128504 199520
rect 127898 192536 127954 192545
rect 127898 192471 127954 192480
rect 127808 180872 127860 180878
rect 127808 180814 127860 180820
rect 127714 179752 127770 179761
rect 127714 179687 127770 179696
rect 127728 179382 127756 179687
rect 127716 179376 127768 179382
rect 127716 179318 127768 179324
rect 127624 155916 127676 155922
rect 127624 155858 127676 155864
rect 126978 148608 127034 148617
rect 126978 148543 127034 148552
rect 127072 146192 127124 146198
rect 127072 146134 127124 146140
rect 126980 144152 127032 144158
rect 126980 144094 127032 144100
rect 126992 143274 127020 144094
rect 126980 143268 127032 143274
rect 126980 143210 127032 143216
rect 126060 142656 126112 142662
rect 126060 142598 126112 142604
rect 126072 139890 126100 142598
rect 127084 139890 127112 146134
rect 127636 143546 127848 143562
rect 127624 143540 127848 143546
rect 127676 143534 127848 143540
rect 127624 143482 127676 143488
rect 127820 143410 127848 143534
rect 127716 143404 127768 143410
rect 127716 143346 127768 143352
rect 127808 143404 127860 143410
rect 127808 143346 127860 143352
rect 127728 139890 127756 143346
rect 126072 139862 126408 139890
rect 127084 139862 127236 139890
rect 127728 139862 128064 139890
rect 128464 139369 128492 199514
rect 128912 198892 128964 198898
rect 128912 198834 128964 198840
rect 128636 194812 128688 194818
rect 128636 194754 128688 194760
rect 128648 192574 128676 194754
rect 128924 193905 128952 198834
rect 129016 197441 129044 200631
rect 177948 200602 178000 200608
rect 132132 200592 132184 200598
rect 132132 200534 132184 200540
rect 131764 200524 131816 200530
rect 131764 200466 131816 200472
rect 131856 200524 131908 200530
rect 131856 200466 131908 200472
rect 131486 200424 131542 200433
rect 131486 200359 131542 200368
rect 131500 200161 131528 200359
rect 131486 200152 131542 200161
rect 131486 200087 131542 200096
rect 131670 200152 131726 200161
rect 131670 200087 131726 200096
rect 129740 200048 129792 200054
rect 129740 199990 129792 199996
rect 129648 199572 129700 199578
rect 129648 199514 129700 199520
rect 129660 199238 129688 199514
rect 129648 199232 129700 199238
rect 129648 199174 129700 199180
rect 129752 198490 129780 199990
rect 131026 199880 131082 199889
rect 131026 199815 131082 199824
rect 130384 199028 130436 199034
rect 130384 198970 130436 198976
rect 129740 198484 129792 198490
rect 129740 198426 129792 198432
rect 129002 197432 129058 197441
rect 129002 197367 129058 197376
rect 128910 193896 128966 193905
rect 128910 193831 128966 193840
rect 128636 192568 128688 192574
rect 128636 192510 128688 192516
rect 128544 142724 128596 142730
rect 128544 142666 128596 142672
rect 128556 139890 128584 142666
rect 128556 139862 128892 139890
rect 124034 139360 124090 139369
rect 124034 139295 124090 139304
rect 125966 139360 126022 139369
rect 125966 139295 126022 139304
rect 128450 139360 128506 139369
rect 129016 139330 129044 197367
rect 129372 146260 129424 146266
rect 129372 146202 129424 146208
rect 129384 139890 129412 146202
rect 130396 146130 130424 198970
rect 131040 197742 131068 199815
rect 131684 199578 131712 200087
rect 131776 199714 131804 200466
rect 131868 200190 131896 200466
rect 132144 200326 132172 200534
rect 177652 200382 177896 200410
rect 132132 200320 132184 200326
rect 132038 200288 132094 200297
rect 132132 200262 132184 200268
rect 132222 200288 132278 200297
rect 132038 200223 132040 200232
rect 132092 200223 132094 200232
rect 132222 200223 132278 200232
rect 132040 200194 132092 200200
rect 131856 200184 131908 200190
rect 131856 200126 131908 200132
rect 131948 200184 132000 200190
rect 131948 200126 132000 200132
rect 131854 200016 131910 200025
rect 131854 199951 131856 199960
rect 131908 199951 131910 199960
rect 131856 199922 131908 199928
rect 131854 199880 131910 199889
rect 131854 199815 131856 199824
rect 131908 199815 131910 199824
rect 131856 199786 131908 199792
rect 131764 199708 131816 199714
rect 131764 199650 131816 199656
rect 131960 199617 131988 200126
rect 132236 199918 132264 200223
rect 177868 200138 177896 200382
rect 177960 200297 177988 200602
rect 178684 200456 178736 200462
rect 178684 200398 178736 200404
rect 178774 200424 178830 200433
rect 177946 200288 178002 200297
rect 177946 200223 178002 200232
rect 132328 200110 132388 200138
rect 132224 199912 132276 199918
rect 132038 199880 132094 199889
rect 132224 199854 132276 199860
rect 132038 199815 132094 199824
rect 131946 199608 132002 199617
rect 131672 199572 131724 199578
rect 131672 199514 131724 199520
rect 131856 199572 131908 199578
rect 131946 199543 132002 199552
rect 131856 199514 131908 199520
rect 131762 197976 131818 197985
rect 131762 197911 131764 197920
rect 131816 197911 131818 197920
rect 131764 197882 131816 197888
rect 131028 197736 131080 197742
rect 131028 197678 131080 197684
rect 131762 197296 131818 197305
rect 131762 197231 131818 197240
rect 130566 195528 130622 195537
rect 130566 195463 130622 195472
rect 130476 190732 130528 190738
rect 130476 190674 130528 190680
rect 130384 146124 130436 146130
rect 130384 146066 130436 146072
rect 130106 146024 130162 146033
rect 130106 145959 130162 145968
rect 130120 139890 130148 145959
rect 130488 140457 130516 190674
rect 130580 144838 130608 195463
rect 130752 195152 130804 195158
rect 130752 195094 130804 195100
rect 130660 194676 130712 194682
rect 130660 194618 130712 194624
rect 130672 148170 130700 194618
rect 130764 148238 130792 195094
rect 130844 186380 130896 186386
rect 130844 186322 130896 186328
rect 130752 148232 130804 148238
rect 130752 148174 130804 148180
rect 130660 148164 130712 148170
rect 130660 148106 130712 148112
rect 130568 144832 130620 144838
rect 130568 144774 130620 144780
rect 130856 141953 130884 186322
rect 131120 177948 131172 177954
rect 131120 177890 131172 177896
rect 131132 177478 131160 177890
rect 131120 177472 131172 177478
rect 131120 177414 131172 177420
rect 131776 148374 131804 197231
rect 131868 197169 131896 199514
rect 131854 197160 131910 197169
rect 131854 197095 131910 197104
rect 131856 196512 131908 196518
rect 131856 196454 131908 196460
rect 131764 148368 131816 148374
rect 131764 148310 131816 148316
rect 131764 146056 131816 146062
rect 131764 145998 131816 146004
rect 131120 142792 131172 142798
rect 131120 142734 131172 142740
rect 131132 142662 131160 142734
rect 131120 142656 131172 142662
rect 131120 142598 131172 142604
rect 130842 141944 130898 141953
rect 130842 141879 130898 141888
rect 130474 140448 130530 140457
rect 130474 140383 130530 140392
rect 131132 139890 131160 142598
rect 131776 139890 131804 145998
rect 131868 140486 131896 196454
rect 131948 196308 132000 196314
rect 131948 196250 132000 196256
rect 131856 140480 131908 140486
rect 131856 140422 131908 140428
rect 131960 140418 131988 196250
rect 132052 194818 132080 199815
rect 132328 197305 132356 200110
rect 132466 199968 132494 200124
rect 132420 199940 132494 199968
rect 132314 197296 132370 197305
rect 132314 197231 132370 197240
rect 132420 197062 132448 199940
rect 132558 199832 132586 200124
rect 132650 199918 132678 200124
rect 132638 199912 132690 199918
rect 132638 199854 132690 199860
rect 132742 199850 132770 200124
rect 132512 199804 132586 199832
rect 132730 199844 132782 199850
rect 132512 198064 132540 199804
rect 132730 199786 132782 199792
rect 132834 199730 132862 200124
rect 132926 199764 132954 200124
rect 133018 199918 133046 200124
rect 133110 199918 133138 200124
rect 133202 199923 133230 200124
rect 133006 199912 133058 199918
rect 133006 199854 133058 199860
rect 133098 199912 133150 199918
rect 133098 199854 133150 199860
rect 133188 199914 133244 199923
rect 133188 199849 133244 199858
rect 133144 199776 133196 199782
rect 132926 199736 133000 199764
rect 132788 199702 132862 199730
rect 132512 198036 132724 198064
rect 132408 197056 132460 197062
rect 132408 196998 132460 197004
rect 132590 196480 132646 196489
rect 132590 196415 132646 196424
rect 132406 196344 132462 196353
rect 132406 196279 132462 196288
rect 132040 194812 132092 194818
rect 132040 194754 132092 194760
rect 132224 194404 132276 194410
rect 132224 194346 132276 194352
rect 132132 188896 132184 188902
rect 132132 188838 132184 188844
rect 132040 187808 132092 187814
rect 132040 187750 132092 187756
rect 132052 140554 132080 187750
rect 132144 140593 132172 188838
rect 132236 148918 132264 194346
rect 132316 193248 132368 193254
rect 132316 193190 132368 193196
rect 132328 193050 132356 193190
rect 132316 193044 132368 193050
rect 132316 192986 132368 192992
rect 132316 192568 132368 192574
rect 132316 192510 132368 192516
rect 132328 148986 132356 192510
rect 132420 177954 132448 196279
rect 132408 177948 132460 177954
rect 132408 177890 132460 177896
rect 132604 151162 132632 196415
rect 132696 191010 132724 198036
rect 132684 191004 132736 191010
rect 132684 190946 132736 190952
rect 132684 190868 132736 190874
rect 132684 190810 132736 190816
rect 132696 151298 132724 190810
rect 132788 177410 132816 199702
rect 132972 192982 133000 199736
rect 133064 199724 133144 199730
rect 133294 199764 133322 200124
rect 133386 199889 133414 200124
rect 133372 199880 133428 199889
rect 133372 199815 133428 199824
rect 133064 199718 133196 199724
rect 133248 199736 133322 199764
rect 133064 199702 133184 199718
rect 132960 192976 133012 192982
rect 132960 192918 133012 192924
rect 132972 192574 133000 192918
rect 132960 192568 133012 192574
rect 132960 192510 133012 192516
rect 132868 191004 132920 191010
rect 132868 190946 132920 190952
rect 132880 178770 132908 190946
rect 133064 180794 133092 199702
rect 133142 199608 133198 199617
rect 133142 199543 133198 199552
rect 133156 198898 133184 199543
rect 133144 198892 133196 198898
rect 133144 198834 133196 198840
rect 133144 197668 133196 197674
rect 133144 197610 133196 197616
rect 132972 180766 133092 180794
rect 132868 178764 132920 178770
rect 132868 178706 132920 178712
rect 132776 177404 132828 177410
rect 132776 177346 132828 177352
rect 132684 151292 132736 151298
rect 132684 151234 132736 151240
rect 132592 151156 132644 151162
rect 132592 151098 132644 151104
rect 132316 148980 132368 148986
rect 132316 148922 132368 148928
rect 132224 148912 132276 148918
rect 132224 148854 132276 148860
rect 132972 148646 133000 180766
rect 132960 148640 133012 148646
rect 132960 148582 133012 148588
rect 132590 145888 132646 145897
rect 132590 145823 132646 145832
rect 132130 140584 132186 140593
rect 132040 140548 132092 140554
rect 132130 140519 132186 140528
rect 132040 140490 132092 140496
rect 131948 140412 132000 140418
rect 131948 140354 132000 140360
rect 132604 139890 132632 145823
rect 133156 140350 133184 197610
rect 133248 195514 133276 199736
rect 133478 199560 133506 200124
rect 133570 199923 133598 200124
rect 133556 199914 133612 199923
rect 133556 199849 133612 199858
rect 133662 199764 133690 200124
rect 133570 199736 133690 199764
rect 133570 199696 133598 199736
rect 133754 199730 133782 200124
rect 133846 199923 133874 200124
rect 133832 199914 133888 199923
rect 133832 199849 133888 199858
rect 133938 199764 133966 200124
rect 134030 199918 134058 200124
rect 134122 199918 134150 200124
rect 134018 199912 134070 199918
rect 134018 199854 134070 199860
rect 134110 199912 134162 199918
rect 134214 199889 134242 200124
rect 134110 199854 134162 199860
rect 134200 199880 134256 199889
rect 134200 199815 134256 199824
rect 134156 199776 134208 199782
rect 133938 199736 134012 199764
rect 133754 199714 133828 199730
rect 133754 199708 133840 199714
rect 133754 199702 133788 199708
rect 133570 199668 133644 199696
rect 133616 199578 133644 199668
rect 133788 199650 133840 199656
rect 133696 199640 133748 199646
rect 133696 199582 133748 199588
rect 133604 199572 133656 199578
rect 133478 199532 133552 199560
rect 133524 198472 133552 199532
rect 133604 199514 133656 199520
rect 133604 199300 133656 199306
rect 133604 199242 133656 199248
rect 133616 199209 133644 199242
rect 133602 199200 133658 199209
rect 133602 199135 133658 199144
rect 133524 198444 133644 198472
rect 133510 198384 133566 198393
rect 133510 198319 133566 198328
rect 133524 197713 133552 198319
rect 133510 197704 133566 197713
rect 133510 197639 133566 197648
rect 133248 195486 133368 195514
rect 133236 195424 133288 195430
rect 133236 195366 133288 195372
rect 133340 195378 133368 195486
rect 133248 194750 133276 195366
rect 133340 195350 133460 195378
rect 133328 195220 133380 195226
rect 133328 195162 133380 195168
rect 133236 194744 133288 194750
rect 133236 194686 133288 194692
rect 133234 190496 133290 190505
rect 133234 190431 133290 190440
rect 133248 190398 133276 190431
rect 133236 190392 133288 190398
rect 133236 190334 133288 190340
rect 133340 180794 133368 195162
rect 133432 194410 133460 195350
rect 133420 194404 133472 194410
rect 133420 194346 133472 194352
rect 133616 193214 133644 198444
rect 133708 198354 133736 199582
rect 133788 199572 133840 199578
rect 133788 199514 133840 199520
rect 133696 198348 133748 198354
rect 133696 198290 133748 198296
rect 133524 193186 133644 193214
rect 133800 193214 133828 199514
rect 133984 197946 134012 199736
rect 134306 199764 134334 200124
rect 134398 199889 134426 200124
rect 134384 199880 134440 199889
rect 134384 199815 134440 199824
rect 134490 199764 134518 200124
rect 134582 199918 134610 200124
rect 134570 199912 134622 199918
rect 134570 199854 134622 199860
rect 134306 199736 134380 199764
rect 134156 199718 134208 199724
rect 134064 199708 134116 199714
rect 134064 199650 134116 199656
rect 134076 199617 134104 199650
rect 134062 199608 134118 199617
rect 134062 199543 134118 199552
rect 133972 197940 134024 197946
rect 133972 197882 134024 197888
rect 133972 197600 134024 197606
rect 133972 197542 134024 197548
rect 133800 193186 133920 193214
rect 133524 191834 133552 193186
rect 133432 191806 133552 191834
rect 133432 190874 133460 191806
rect 133892 191418 133920 193186
rect 133880 191412 133932 191418
rect 133880 191354 133932 191360
rect 133420 190868 133472 190874
rect 133420 190810 133472 190816
rect 133984 189990 134012 197542
rect 134168 191834 134196 199718
rect 134352 199578 134380 199736
rect 134444 199736 134518 199764
rect 134674 199764 134702 200124
rect 134766 199889 134794 200124
rect 134752 199880 134808 199889
rect 134752 199815 134808 199824
rect 134858 199764 134886 200124
rect 134950 199918 134978 200124
rect 134938 199912 134990 199918
rect 134938 199854 134990 199860
rect 134674 199736 134748 199764
rect 134340 199572 134392 199578
rect 134340 199514 134392 199520
rect 134444 198286 134472 199736
rect 134524 199640 134576 199646
rect 134524 199582 134576 199588
rect 134536 198694 134564 199582
rect 134524 198688 134576 198694
rect 134524 198630 134576 198636
rect 134616 198484 134668 198490
rect 134616 198426 134668 198432
rect 134432 198280 134484 198286
rect 134628 198257 134656 198426
rect 134432 198222 134484 198228
rect 134614 198248 134670 198257
rect 134614 198183 134670 198192
rect 134432 195968 134484 195974
rect 134432 195910 134484 195916
rect 134338 193352 134394 193361
rect 134338 193287 134394 193296
rect 134168 191806 134288 191834
rect 134064 191004 134116 191010
rect 134064 190946 134116 190952
rect 133972 189984 134024 189990
rect 133972 189926 134024 189932
rect 133248 180766 133368 180794
rect 133248 148850 133276 180766
rect 133788 179308 133840 179314
rect 133788 179250 133840 179256
rect 133800 178770 133828 179250
rect 133788 178764 133840 178770
rect 133788 178706 133840 178712
rect 133788 178016 133840 178022
rect 133788 177958 133840 177964
rect 133800 177410 133828 177958
rect 133788 177404 133840 177410
rect 133788 177346 133840 177352
rect 134076 151094 134104 190946
rect 134064 151088 134116 151094
rect 134064 151030 134116 151036
rect 133236 148844 133288 148850
rect 133236 148786 133288 148792
rect 134260 148714 134288 191806
rect 134352 151230 134380 193287
rect 134444 191758 134472 195910
rect 134720 194313 134748 199736
rect 134812 199736 134886 199764
rect 134706 194304 134762 194313
rect 134706 194239 134762 194248
rect 134524 193248 134576 193254
rect 134524 193190 134576 193196
rect 134432 191752 134484 191758
rect 134432 191694 134484 191700
rect 134340 151224 134392 151230
rect 134340 151166 134392 151172
rect 134248 148708 134300 148714
rect 134248 148650 134300 148656
rect 134248 145988 134300 145994
rect 134248 145930 134300 145936
rect 133512 143472 133564 143478
rect 133512 143414 133564 143420
rect 133144 140344 133196 140350
rect 133144 140286 133196 140292
rect 133524 139890 133552 143414
rect 134260 139890 134288 145930
rect 134536 141817 134564 193190
rect 134812 191010 134840 199736
rect 134892 199640 134944 199646
rect 135042 199628 135070 200124
rect 135134 199923 135162 200124
rect 135120 199914 135176 199923
rect 135120 199849 135176 199858
rect 135226 199764 135254 200124
rect 134892 199582 134944 199588
rect 134996 199600 135070 199628
rect 135180 199736 135254 199764
rect 134904 195673 134932 199582
rect 134890 195664 134946 195673
rect 134890 195599 134946 195608
rect 134800 191004 134852 191010
rect 134800 190946 134852 190952
rect 134996 187066 135024 199600
rect 135076 199300 135128 199306
rect 135076 199242 135128 199248
rect 135088 196761 135116 199242
rect 135074 196752 135130 196761
rect 135074 196687 135130 196696
rect 135180 195974 135208 199736
rect 135318 199696 135346 200124
rect 135410 199918 135438 200124
rect 135398 199912 135450 199918
rect 135502 199889 135530 200124
rect 135398 199854 135450 199860
rect 135488 199880 135544 199889
rect 135488 199815 135544 199824
rect 135594 199764 135622 200124
rect 135686 199889 135714 200124
rect 135778 199918 135806 200124
rect 135766 199912 135818 199918
rect 135672 199880 135728 199889
rect 135766 199854 135818 199860
rect 135672 199815 135728 199824
rect 135870 199764 135898 200124
rect 135272 199668 135346 199696
rect 135442 199744 135498 199753
rect 135594 199736 135668 199764
rect 135442 199679 135498 199688
rect 135272 197985 135300 199668
rect 135352 199572 135404 199578
rect 135352 199514 135404 199520
rect 135258 197976 135314 197985
rect 135258 197911 135314 197920
rect 135168 195968 135220 195974
rect 135168 195910 135220 195916
rect 135364 191834 135392 199514
rect 135456 192710 135484 199679
rect 135534 199608 135590 199617
rect 135534 199543 135590 199552
rect 135548 195498 135576 199543
rect 135640 199306 135668 199736
rect 135824 199736 135898 199764
rect 135962 199753 135990 200124
rect 136054 199918 136082 200124
rect 136146 199918 136174 200124
rect 136238 199918 136266 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136134 199912 136186 199918
rect 136134 199854 136186 199860
rect 136226 199912 136278 199918
rect 136226 199854 136278 199860
rect 136088 199776 136140 199782
rect 135948 199744 136004 199753
rect 135720 199640 135772 199646
rect 135720 199582 135772 199588
rect 135628 199300 135680 199306
rect 135628 199242 135680 199248
rect 135536 195492 135588 195498
rect 135536 195434 135588 195440
rect 135444 192704 135496 192710
rect 135444 192646 135496 192652
rect 135732 191834 135760 199582
rect 135824 193730 135852 199736
rect 136088 199718 136140 199724
rect 136180 199776 136232 199782
rect 136330 199764 136358 200124
rect 136422 199918 136450 200124
rect 136410 199912 136462 199918
rect 136514 199889 136542 200124
rect 136410 199854 136462 199860
rect 136500 199880 136556 199889
rect 136500 199815 136556 199824
rect 136606 199764 136634 200124
rect 136698 199850 136726 200124
rect 136686 199844 136738 199850
rect 136686 199786 136738 199792
rect 136180 199718 136232 199724
rect 136284 199736 136358 199764
rect 136560 199736 136634 199764
rect 135948 199679 136004 199688
rect 135996 199096 136048 199102
rect 135996 199038 136048 199044
rect 135904 198892 135956 198898
rect 135904 198834 135956 198840
rect 135916 198801 135944 198834
rect 135902 198792 135958 198801
rect 135902 198727 135958 198736
rect 136008 198082 136036 199038
rect 135996 198076 136048 198082
rect 135996 198018 136048 198024
rect 135904 197056 135956 197062
rect 135904 196998 135956 197004
rect 135812 193724 135864 193730
rect 135812 193666 135864 193672
rect 135364 191806 135668 191834
rect 135732 191806 135852 191834
rect 135536 191412 135588 191418
rect 135536 191354 135588 191360
rect 134984 187060 135036 187066
rect 134984 187002 135036 187008
rect 135548 184006 135576 191354
rect 135536 184000 135588 184006
rect 135536 183942 135588 183948
rect 135640 147014 135668 191806
rect 135720 191004 135772 191010
rect 135720 190946 135772 190952
rect 135732 148510 135760 190946
rect 135824 187066 135852 191806
rect 135812 187060 135864 187066
rect 135812 187002 135864 187008
rect 135916 184142 135944 196998
rect 136100 191834 136128 199718
rect 136192 195945 136220 199718
rect 136284 199209 136312 199736
rect 136456 199708 136508 199714
rect 136456 199650 136508 199656
rect 136364 199640 136416 199646
rect 136364 199582 136416 199588
rect 136270 199200 136326 199209
rect 136270 199135 136326 199144
rect 136272 198688 136324 198694
rect 136272 198630 136324 198636
rect 136178 195936 136234 195945
rect 136178 195871 136234 195880
rect 136100 191806 136220 191834
rect 136192 187542 136220 191806
rect 136284 190058 136312 198630
rect 136376 197062 136404 199582
rect 136468 197062 136496 199650
rect 136364 197056 136416 197062
rect 136364 196998 136416 197004
rect 136456 197056 136508 197062
rect 136456 196998 136508 197004
rect 136364 196716 136416 196722
rect 136364 196658 136416 196664
rect 136376 192642 136404 196658
rect 136454 195936 136510 195945
rect 136454 195871 136510 195880
rect 136364 192636 136416 192642
rect 136364 192578 136416 192584
rect 136468 191010 136496 195871
rect 136560 191418 136588 199736
rect 136790 199730 136818 200124
rect 136882 199889 136910 200124
rect 136868 199880 136924 199889
rect 136868 199815 136924 199824
rect 136744 199702 136818 199730
rect 136638 198248 136694 198257
rect 136638 198183 136694 198192
rect 136652 197849 136680 198183
rect 136638 197840 136694 197849
rect 136638 197775 136694 197784
rect 136640 197056 136692 197062
rect 136640 196998 136692 197004
rect 136652 196722 136680 196998
rect 136640 196716 136692 196722
rect 136640 196658 136692 196664
rect 136638 196072 136694 196081
rect 136638 196007 136694 196016
rect 136652 195401 136680 196007
rect 136744 195945 136772 199702
rect 136974 199628 137002 200124
rect 137066 199730 137094 200124
rect 137158 199850 137186 200124
rect 137250 199918 137278 200124
rect 137238 199912 137290 199918
rect 137238 199854 137290 199860
rect 137342 199850 137370 200124
rect 137146 199844 137198 199850
rect 137146 199786 137198 199792
rect 137330 199844 137382 199850
rect 137330 199786 137382 199792
rect 137434 199730 137462 200124
rect 137066 199702 137140 199730
rect 136822 199608 136878 199617
rect 136822 199543 136878 199552
rect 136928 199600 137002 199628
rect 136836 198422 136864 199543
rect 136824 198416 136876 198422
rect 136824 198358 136876 198364
rect 136822 197840 136878 197849
rect 136822 197775 136878 197784
rect 136836 197441 136864 197775
rect 136822 197432 136878 197441
rect 136822 197367 136878 197376
rect 136730 195936 136786 195945
rect 136730 195871 136786 195880
rect 136638 195392 136694 195401
rect 136638 195327 136694 195336
rect 136928 191826 136956 199600
rect 137112 199424 137140 199702
rect 137192 199708 137244 199714
rect 137192 199650 137244 199656
rect 137284 199708 137336 199714
rect 137284 199650 137336 199656
rect 137388 199702 137462 199730
rect 137526 199730 137554 200124
rect 137618 199918 137646 200124
rect 137710 199918 137738 200124
rect 137802 199918 137830 200124
rect 137606 199912 137658 199918
rect 137606 199854 137658 199860
rect 137698 199912 137750 199918
rect 137698 199854 137750 199860
rect 137790 199912 137842 199918
rect 137894 199889 137922 200124
rect 137986 199918 138014 200124
rect 137974 199912 138026 199918
rect 137790 199854 137842 199860
rect 137880 199880 137936 199889
rect 137974 199854 138026 199860
rect 137880 199815 137936 199824
rect 137652 199776 137704 199782
rect 137526 199702 137600 199730
rect 137652 199718 137704 199724
rect 137020 199396 137140 199424
rect 136916 191820 136968 191826
rect 136916 191762 136968 191768
rect 136548 191412 136600 191418
rect 136548 191354 136600 191360
rect 137020 191162 137048 199396
rect 137098 198656 137154 198665
rect 137098 198591 137154 198600
rect 137112 193934 137140 198591
rect 137204 198529 137232 199650
rect 137190 198520 137246 198529
rect 137190 198455 137246 198464
rect 137192 196104 137244 196110
rect 137192 196046 137244 196052
rect 137100 193928 137152 193934
rect 137100 193870 137152 193876
rect 137204 191758 137232 196046
rect 137296 195974 137324 199650
rect 137388 196217 137416 199702
rect 137468 199572 137520 199578
rect 137468 199514 137520 199520
rect 137374 196208 137430 196217
rect 137374 196143 137430 196152
rect 137480 196110 137508 199514
rect 137468 196104 137520 196110
rect 137468 196046 137520 196052
rect 137296 195946 137508 195974
rect 137376 195492 137428 195498
rect 137376 195434 137428 195440
rect 137192 191752 137244 191758
rect 137192 191694 137244 191700
rect 137100 191412 137152 191418
rect 137100 191354 137152 191360
rect 136836 191134 137048 191162
rect 136456 191004 136508 191010
rect 136456 190946 136508 190952
rect 136640 190460 136692 190466
rect 136640 190402 136692 190408
rect 136272 190052 136324 190058
rect 136272 189994 136324 190000
rect 136652 189174 136680 190402
rect 136640 189168 136692 189174
rect 136640 189110 136692 189116
rect 136180 187536 136232 187542
rect 136180 187478 136232 187484
rect 136180 187060 136232 187066
rect 136180 187002 136232 187008
rect 135904 184136 135956 184142
rect 135904 184078 135956 184084
rect 136192 180674 136220 187002
rect 136180 180668 136232 180674
rect 136180 180610 136232 180616
rect 136192 180334 136220 180610
rect 136180 180328 136232 180334
rect 136180 180270 136232 180276
rect 136546 179480 136602 179489
rect 136546 179415 136602 179424
rect 136454 177848 136510 177857
rect 136560 177818 136588 179415
rect 136454 177783 136510 177792
rect 136548 177812 136600 177818
rect 136468 176662 136496 177783
rect 136548 177754 136600 177760
rect 136560 177342 136588 177754
rect 136548 177336 136600 177342
rect 136548 177278 136600 177284
rect 136456 176656 136508 176662
rect 136456 176598 136508 176604
rect 136468 175982 136496 176598
rect 136836 176225 136864 191134
rect 137008 190868 137060 190874
rect 137008 190810 137060 190816
rect 136916 190800 136968 190806
rect 136916 190742 136968 190748
rect 136928 180470 136956 190742
rect 137020 180606 137048 190810
rect 137112 181762 137140 191354
rect 137388 190806 137416 195434
rect 137376 190800 137428 190806
rect 137376 190742 137428 190748
rect 137192 190664 137244 190670
rect 137192 190606 137244 190612
rect 137100 181756 137152 181762
rect 137100 181698 137152 181704
rect 137008 180600 137060 180606
rect 137008 180542 137060 180548
rect 136916 180464 136968 180470
rect 136916 180406 136968 180412
rect 136928 180130 136956 180406
rect 137020 180198 137048 180542
rect 137008 180192 137060 180198
rect 137008 180134 137060 180140
rect 136916 180124 136968 180130
rect 136916 180066 136968 180072
rect 136822 176216 136878 176225
rect 136822 176151 136878 176160
rect 136456 175976 136508 175982
rect 136456 175918 136508 175924
rect 135720 148504 135772 148510
rect 135720 148446 135772 148452
rect 135628 147008 135680 147014
rect 135628 146950 135680 146956
rect 135260 145920 135312 145926
rect 135260 145862 135312 145868
rect 134522 141808 134578 141817
rect 134522 141743 134578 141752
rect 135272 139890 135300 145862
rect 136730 145752 136786 145761
rect 136730 145687 136786 145696
rect 135994 143032 136050 143041
rect 135994 142967 136050 142976
rect 136008 139890 136036 142967
rect 136744 139890 136772 145687
rect 137204 140146 137232 190606
rect 137284 190460 137336 190466
rect 137284 190402 137336 190408
rect 137296 190369 137324 190402
rect 137282 190360 137338 190369
rect 137282 190295 137338 190304
rect 137282 179480 137338 179489
rect 137282 179415 137338 179424
rect 137296 140729 137324 179415
rect 137480 146946 137508 195946
rect 137572 190874 137600 199702
rect 137664 195498 137692 199718
rect 137744 199708 137796 199714
rect 137744 199650 137796 199656
rect 137652 195492 137704 195498
rect 137652 195434 137704 195440
rect 137652 191820 137704 191826
rect 137652 191762 137704 191768
rect 137560 190868 137612 190874
rect 137560 190810 137612 190816
rect 137664 186314 137692 191762
rect 137756 191418 137784 199650
rect 137836 199640 137888 199646
rect 138078 199628 138106 200124
rect 138170 199889 138198 200124
rect 138156 199880 138212 199889
rect 138156 199815 138212 199824
rect 138262 199696 138290 200124
rect 138354 199764 138382 200124
rect 138446 199889 138474 200124
rect 138432 199880 138488 199889
rect 138432 199815 138488 199824
rect 138354 199736 138428 199764
rect 137836 199582 137888 199588
rect 137926 199608 137982 199617
rect 137848 199209 137876 199582
rect 137926 199543 137982 199552
rect 138032 199600 138106 199628
rect 138216 199668 138290 199696
rect 137834 199200 137890 199209
rect 137834 199135 137890 199144
rect 137940 198880 137968 199543
rect 138032 199306 138060 199600
rect 138020 199300 138072 199306
rect 138020 199242 138072 199248
rect 137848 198852 137968 198880
rect 137744 191412 137796 191418
rect 137744 191354 137796 191360
rect 137848 190670 137876 198852
rect 138032 198778 138060 199242
rect 137940 198750 138060 198778
rect 137940 195226 137968 198750
rect 138018 198520 138074 198529
rect 138018 198455 138074 198464
rect 138032 198014 138060 198455
rect 138020 198008 138072 198014
rect 138020 197950 138072 197956
rect 138216 197810 138244 199668
rect 138296 199572 138348 199578
rect 138296 199514 138348 199520
rect 138308 198336 138336 199514
rect 138400 198626 138428 199736
rect 138538 199696 138566 200124
rect 138630 199764 138658 200124
rect 138722 199918 138750 200124
rect 138814 199918 138842 200124
rect 138906 199918 138934 200124
rect 138710 199912 138762 199918
rect 138710 199854 138762 199860
rect 138802 199912 138854 199918
rect 138802 199854 138854 199860
rect 138894 199912 138946 199918
rect 138894 199854 138946 199860
rect 138848 199776 138900 199782
rect 138630 199736 138704 199764
rect 138538 199668 138612 199696
rect 138480 199572 138532 199578
rect 138480 199514 138532 199520
rect 138388 198620 138440 198626
rect 138388 198562 138440 198568
rect 138308 198308 138428 198336
rect 138294 198248 138350 198257
rect 138294 198183 138350 198192
rect 138204 197804 138256 197810
rect 138204 197746 138256 197752
rect 138308 197577 138336 198183
rect 138294 197568 138350 197577
rect 138020 197532 138072 197538
rect 138294 197503 138350 197512
rect 138020 197474 138072 197480
rect 137928 195220 137980 195226
rect 137928 195162 137980 195168
rect 138032 193118 138060 197474
rect 138202 196752 138258 196761
rect 138202 196687 138258 196696
rect 138112 196104 138164 196110
rect 138112 196046 138164 196052
rect 138020 193112 138072 193118
rect 138020 193054 138072 193060
rect 137928 191752 137980 191758
rect 137928 191694 137980 191700
rect 137836 190664 137888 190670
rect 137836 190606 137888 190612
rect 137572 186286 137692 186314
rect 137572 181626 137600 186286
rect 137940 181694 137968 191694
rect 138124 190454 138152 196046
rect 138216 192846 138244 196687
rect 138400 196217 138428 198308
rect 138386 196208 138442 196217
rect 138492 196178 138520 199514
rect 138584 196926 138612 199668
rect 138572 196920 138624 196926
rect 138572 196862 138624 196868
rect 138386 196143 138442 196152
rect 138480 196172 138532 196178
rect 138480 196114 138532 196120
rect 138676 196058 138704 199736
rect 138768 199736 138848 199764
rect 138768 198257 138796 199736
rect 138848 199718 138900 199724
rect 138998 199696 139026 200124
rect 139090 199889 139118 200124
rect 139182 199918 139210 200124
rect 139170 199912 139222 199918
rect 139076 199880 139132 199889
rect 139170 199854 139222 199860
rect 139076 199815 139132 199824
rect 139274 199764 139302 200124
rect 139366 199889 139394 200124
rect 139458 199918 139486 200124
rect 139446 199912 139498 199918
rect 139352 199880 139408 199889
rect 139550 199889 139578 200124
rect 139446 199854 139498 199860
rect 139536 199880 139592 199889
rect 139352 199815 139408 199824
rect 139536 199815 139592 199824
rect 139228 199736 139302 199764
rect 139400 199776 139452 199782
rect 138998 199668 139072 199696
rect 138848 199572 138900 199578
rect 138848 199514 138900 199520
rect 138754 198248 138810 198257
rect 138754 198183 138810 198192
rect 138756 197872 138808 197878
rect 138756 197814 138808 197820
rect 138768 197538 138796 197814
rect 138756 197532 138808 197538
rect 138756 197474 138808 197480
rect 138756 196784 138808 196790
rect 138756 196726 138808 196732
rect 138308 196030 138704 196058
rect 138204 192840 138256 192846
rect 138204 192782 138256 192788
rect 138032 190426 138152 190454
rect 138032 186250 138060 190426
rect 138020 186244 138072 186250
rect 138020 186186 138072 186192
rect 138032 185638 138060 186186
rect 138308 185706 138336 196030
rect 138480 195968 138532 195974
rect 138386 195936 138442 195945
rect 138480 195910 138532 195916
rect 138386 195871 138442 195880
rect 138296 185700 138348 185706
rect 138296 185642 138348 185648
rect 138020 185632 138072 185638
rect 138020 185574 138072 185580
rect 137928 181688 137980 181694
rect 137928 181630 137980 181636
rect 137560 181620 137612 181626
rect 137560 181562 137612 181568
rect 137468 146940 137520 146946
rect 137468 146882 137520 146888
rect 137928 144220 137980 144226
rect 137928 144162 137980 144168
rect 137282 140720 137338 140729
rect 137282 140655 137338 140664
rect 137192 140140 137244 140146
rect 137192 140082 137244 140088
rect 137940 139890 137968 144162
rect 138400 140078 138428 195871
rect 138492 141914 138520 195910
rect 138768 191834 138796 196726
rect 138676 191806 138796 191834
rect 138676 144906 138704 191806
rect 138860 180794 138888 199514
rect 138940 199504 138992 199510
rect 138940 199446 138992 199452
rect 138952 199102 138980 199446
rect 138940 199096 138992 199102
rect 139044 199073 139072 199668
rect 139124 199640 139176 199646
rect 139124 199582 139176 199588
rect 138940 199038 138992 199044
rect 139030 199064 139086 199073
rect 139030 198999 139086 199008
rect 138938 197432 138994 197441
rect 138938 197367 138994 197376
rect 138952 196314 138980 197367
rect 138940 196308 138992 196314
rect 138940 196250 138992 196256
rect 139136 195945 139164 199582
rect 139122 195936 139178 195945
rect 139122 195871 139178 195880
rect 139030 183560 139086 183569
rect 139030 183495 139086 183504
rect 138768 180766 138888 180794
rect 138768 179246 138796 180766
rect 138756 179240 138808 179246
rect 138756 179182 138808 179188
rect 138768 178702 138796 179182
rect 139044 179178 139072 183495
rect 139228 182850 139256 199736
rect 139642 199764 139670 200124
rect 139734 199918 139762 200124
rect 139722 199912 139774 199918
rect 139722 199854 139774 199860
rect 139826 199764 139854 200124
rect 139918 199918 139946 200124
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 140010 199764 140038 200124
rect 140102 199889 140130 200124
rect 140088 199880 140144 199889
rect 140088 199815 140144 199824
rect 139400 199718 139452 199724
rect 139596 199736 139670 199764
rect 139780 199736 139854 199764
rect 139964 199736 140038 199764
rect 140194 199764 140222 200124
rect 140286 199889 140314 200124
rect 140272 199880 140328 199889
rect 140272 199815 140328 199824
rect 140378 199764 140406 200124
rect 140470 199918 140498 200124
rect 140458 199912 140510 199918
rect 140458 199854 140510 199860
rect 140562 199764 140590 200124
rect 140654 199918 140682 200124
rect 140642 199912 140694 199918
rect 140642 199854 140694 199860
rect 140746 199764 140774 200124
rect 140838 199918 140866 200124
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140930 199764 140958 200124
rect 140194 199753 140268 199764
rect 140194 199744 140282 199753
rect 140194 199736 140226 199744
rect 139306 199200 139362 199209
rect 139306 199135 139362 199144
rect 139320 191834 139348 199135
rect 139412 195498 139440 199718
rect 139492 199640 139544 199646
rect 139492 199582 139544 199588
rect 139504 197520 139532 199582
rect 139596 197946 139624 199736
rect 139676 199640 139728 199646
rect 139676 199582 139728 199588
rect 139688 198121 139716 199582
rect 139674 198112 139730 198121
rect 139674 198047 139730 198056
rect 139584 197940 139636 197946
rect 139584 197882 139636 197888
rect 139504 197492 139716 197520
rect 139492 197396 139544 197402
rect 139492 197338 139544 197344
rect 139400 195492 139452 195498
rect 139400 195434 139452 195440
rect 139504 195158 139532 197338
rect 139584 196716 139636 196722
rect 139584 196658 139636 196664
rect 139492 195152 139544 195158
rect 139492 195094 139544 195100
rect 139320 191806 139532 191834
rect 139400 191752 139452 191758
rect 139400 191694 139452 191700
rect 139412 191146 139440 191694
rect 139400 191140 139452 191146
rect 139400 191082 139452 191088
rect 139504 189786 139532 191806
rect 139492 189780 139544 189786
rect 139492 189722 139544 189728
rect 139596 184074 139624 196658
rect 139688 184414 139716 197492
rect 139780 192438 139808 199736
rect 139860 199640 139912 199646
rect 139860 199582 139912 199588
rect 139768 192432 139820 192438
rect 139768 192374 139820 192380
rect 139872 189038 139900 199582
rect 139964 196110 139992 199736
rect 140378 199736 140452 199764
rect 140226 199679 140282 199688
rect 140320 199640 140372 199646
rect 140042 199608 140098 199617
rect 140320 199582 140372 199588
rect 140042 199543 140098 199552
rect 140056 199374 140084 199543
rect 140044 199368 140096 199374
rect 140044 199310 140096 199316
rect 140042 199200 140098 199209
rect 140042 199135 140098 199144
rect 140056 197656 140084 199135
rect 140056 197628 140176 197656
rect 140044 197532 140096 197538
rect 140044 197474 140096 197480
rect 139952 196104 140004 196110
rect 139952 196046 140004 196052
rect 139952 195968 140004 195974
rect 139952 195910 140004 195916
rect 139860 189032 139912 189038
rect 139860 188974 139912 188980
rect 139676 184408 139728 184414
rect 139676 184350 139728 184356
rect 139584 184068 139636 184074
rect 139584 184010 139636 184016
rect 139216 182844 139268 182850
rect 139216 182786 139268 182792
rect 139032 179172 139084 179178
rect 139032 179114 139084 179120
rect 138756 178696 138808 178702
rect 138756 178638 138808 178644
rect 138664 144900 138716 144906
rect 138664 144842 138716 144848
rect 138572 143404 138624 143410
rect 138572 143346 138624 143352
rect 138480 141908 138532 141914
rect 138480 141850 138532 141856
rect 138388 140072 138440 140078
rect 138388 140014 138440 140020
rect 138584 139890 138612 143346
rect 139400 143336 139452 143342
rect 139400 143278 139452 143284
rect 139412 139890 139440 143278
rect 139964 141574 139992 195910
rect 140056 194682 140084 197474
rect 140044 194676 140096 194682
rect 140044 194618 140096 194624
rect 140044 193112 140096 193118
rect 140044 193054 140096 193060
rect 140056 192234 140084 193054
rect 140044 192228 140096 192234
rect 140044 192170 140096 192176
rect 140148 190454 140176 197628
rect 140332 196314 140360 199582
rect 140320 196308 140372 196314
rect 140320 196250 140372 196256
rect 140424 195974 140452 199736
rect 140516 199736 140590 199764
rect 140700 199736 140774 199764
rect 140884 199736 140958 199764
rect 141022 199764 141050 200124
rect 141114 199918 141142 200124
rect 141206 199918 141234 200124
rect 141298 199918 141326 200124
rect 141390 199918 141418 200124
rect 141102 199912 141154 199918
rect 141102 199854 141154 199860
rect 141194 199912 141246 199918
rect 141194 199854 141246 199860
rect 141286 199912 141338 199918
rect 141286 199854 141338 199860
rect 141378 199912 141430 199918
rect 141482 199889 141510 200124
rect 141378 199854 141430 199860
rect 141468 199880 141524 199889
rect 141468 199815 141524 199824
rect 141240 199776 141292 199782
rect 141022 199736 141096 199764
rect 140516 196761 140544 199736
rect 140596 199436 140648 199442
rect 140596 199378 140648 199384
rect 140502 196752 140558 196761
rect 140502 196687 140558 196696
rect 140412 195968 140464 195974
rect 140412 195910 140464 195916
rect 140412 195492 140464 195498
rect 140412 195434 140464 195440
rect 140148 190426 140360 190454
rect 140332 147082 140360 190426
rect 140424 185570 140452 195434
rect 140608 191834 140636 199378
rect 140700 196722 140728 199736
rect 140780 199436 140832 199442
rect 140780 199378 140832 199384
rect 140688 196716 140740 196722
rect 140688 196658 140740 196664
rect 140792 196518 140820 199378
rect 140884 198490 140912 199736
rect 141068 199646 141096 199736
rect 141240 199718 141292 199724
rect 141574 199730 141602 200124
rect 141666 199889 141694 200124
rect 141652 199880 141708 199889
rect 141652 199815 141708 199824
rect 141148 199708 141200 199714
rect 141148 199650 141200 199656
rect 140964 199640 141016 199646
rect 140964 199582 141016 199588
rect 141056 199640 141108 199646
rect 141056 199582 141108 199588
rect 140976 198898 141004 199582
rect 141056 199504 141108 199510
rect 141056 199446 141108 199452
rect 140964 198892 141016 198898
rect 140964 198834 141016 198840
rect 140872 198484 140924 198490
rect 140872 198426 140924 198432
rect 140962 198248 141018 198257
rect 140962 198183 141018 198192
rect 140870 197840 140926 197849
rect 140870 197775 140926 197784
rect 140780 196512 140832 196518
rect 140780 196454 140832 196460
rect 140608 191806 140728 191834
rect 140700 191758 140728 191806
rect 140688 191752 140740 191758
rect 140688 191694 140740 191700
rect 140412 185564 140464 185570
rect 140412 185506 140464 185512
rect 140780 176588 140832 176594
rect 140780 176530 140832 176536
rect 140792 176050 140820 176530
rect 140884 176089 140912 197775
rect 140976 196602 141004 198183
rect 141068 196790 141096 199446
rect 141056 196784 141108 196790
rect 141056 196726 141108 196732
rect 140976 196574 141096 196602
rect 140964 195152 141016 195158
rect 140964 195094 141016 195100
rect 140976 176497 141004 195094
rect 141068 176594 141096 196574
rect 141160 194970 141188 199650
rect 141252 196489 141280 199718
rect 141332 199708 141384 199714
rect 141574 199702 141648 199730
rect 141332 199650 141384 199656
rect 141238 196480 141294 196489
rect 141238 196415 141294 196424
rect 141344 195158 141372 199650
rect 141516 199640 141568 199646
rect 141516 199582 141568 199588
rect 141424 199232 141476 199238
rect 141424 199174 141476 199180
rect 141436 198801 141464 199174
rect 141422 198792 141478 198801
rect 141422 198727 141478 198736
rect 141528 198422 141556 199582
rect 141516 198416 141568 198422
rect 141516 198358 141568 198364
rect 141424 197736 141476 197742
rect 141424 197678 141476 197684
rect 141332 195152 141384 195158
rect 141332 195094 141384 195100
rect 141160 194942 141280 194970
rect 141148 194880 141200 194886
rect 141148 194822 141200 194828
rect 141160 183394 141188 194822
rect 141252 194750 141280 194942
rect 141240 194744 141292 194750
rect 141240 194686 141292 194692
rect 141436 190454 141464 197678
rect 141620 196450 141648 199702
rect 141758 199696 141786 200124
rect 141850 199730 141878 200124
rect 141942 199918 141970 200124
rect 141930 199912 141982 199918
rect 141930 199854 141982 199860
rect 142034 199764 142062 200124
rect 142126 199889 142154 200124
rect 142218 199918 142246 200124
rect 142310 199918 142338 200124
rect 142402 199918 142430 200124
rect 142206 199912 142258 199918
rect 142112 199880 142168 199889
rect 142206 199854 142258 199860
rect 142298 199912 142350 199918
rect 142298 199854 142350 199860
rect 142390 199912 142442 199918
rect 142494 199889 142522 200124
rect 142586 199918 142614 200124
rect 142678 199918 142706 200124
rect 142770 199918 142798 200124
rect 142862 199918 142890 200124
rect 142574 199912 142626 199918
rect 142390 199854 142442 199860
rect 142480 199880 142536 199889
rect 142112 199815 142168 199824
rect 142574 199854 142626 199860
rect 142666 199912 142718 199918
rect 142666 199854 142718 199860
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142850 199912 142902 199918
rect 142954 199889 142982 200124
rect 142850 199854 142902 199860
rect 142940 199880 142996 199889
rect 142480 199815 142536 199824
rect 142940 199815 142996 199824
rect 141988 199736 142062 199764
rect 142160 199776 142212 199782
rect 141850 199702 141924 199730
rect 141712 199668 141786 199696
rect 141608 196444 141660 196450
rect 141608 196386 141660 196392
rect 141608 196308 141660 196314
rect 141608 196250 141660 196256
rect 141516 191820 141568 191826
rect 141516 191762 141568 191768
rect 141528 190738 141556 191762
rect 141516 190732 141568 190738
rect 141516 190674 141568 190680
rect 141620 190454 141648 196250
rect 141712 194886 141740 199668
rect 141896 194886 141924 199702
rect 141988 197169 142016 199736
rect 142436 199776 142488 199782
rect 142160 199718 142212 199724
rect 142434 199744 142436 199753
rect 142620 199776 142672 199782
rect 142488 199744 142490 199753
rect 142172 198393 142200 199718
rect 142252 199708 142304 199714
rect 142620 199718 142672 199724
rect 142896 199776 142948 199782
rect 143046 199764 143074 200124
rect 142896 199718 142948 199724
rect 143000 199736 143074 199764
rect 143138 199764 143166 200124
rect 143230 199889 143258 200124
rect 143216 199880 143272 199889
rect 143216 199815 143272 199824
rect 143322 199764 143350 200124
rect 143138 199736 143212 199764
rect 143276 199753 143350 199764
rect 142434 199679 142490 199688
rect 142528 199708 142580 199714
rect 142252 199650 142304 199656
rect 142528 199650 142580 199656
rect 142264 198529 142292 199650
rect 142342 199608 142398 199617
rect 142342 199543 142398 199552
rect 142436 199572 142488 199578
rect 142250 198520 142306 198529
rect 142250 198455 142306 198464
rect 142158 198384 142214 198393
rect 142158 198319 142214 198328
rect 142356 198234 142384 199543
rect 142436 199514 142488 199520
rect 142448 198490 142476 199514
rect 142436 198484 142488 198490
rect 142436 198426 142488 198432
rect 142080 198206 142384 198234
rect 141974 197160 142030 197169
rect 141974 197095 142030 197104
rect 141976 196716 142028 196722
rect 141976 196658 142028 196664
rect 141700 194880 141752 194886
rect 141700 194822 141752 194828
rect 141884 194880 141936 194886
rect 141884 194822 141936 194828
rect 141988 193214 142016 196658
rect 142080 193798 142108 198206
rect 142252 198144 142304 198150
rect 142252 198086 142304 198092
rect 142160 196580 142212 196586
rect 142160 196522 142212 196528
rect 142068 193792 142120 193798
rect 142068 193734 142120 193740
rect 141988 193186 142108 193214
rect 142172 193186 142200 196522
rect 141436 190426 141556 190454
rect 141620 190426 141740 190454
rect 141148 183388 141200 183394
rect 141148 183330 141200 183336
rect 141422 177984 141478 177993
rect 141422 177919 141478 177928
rect 141056 176588 141108 176594
rect 141056 176530 141108 176536
rect 140962 176488 141018 176497
rect 140962 176423 141018 176432
rect 140870 176080 140926 176089
rect 140780 176044 140832 176050
rect 140870 176015 140926 176024
rect 140780 175986 140832 175992
rect 140320 147076 140372 147082
rect 140320 147018 140372 147024
rect 140136 144764 140188 144770
rect 140136 144706 140188 144712
rect 139952 141568 140004 141574
rect 139952 141510 140004 141516
rect 140148 139890 140176 144706
rect 140964 143200 141016 143206
rect 140964 143142 141016 143148
rect 140976 139890 141004 143142
rect 129384 139862 129720 139890
rect 130120 139862 130548 139890
rect 131132 139862 131376 139890
rect 131776 139862 132204 139890
rect 132604 139862 133032 139890
rect 133524 139862 133860 139890
rect 134260 139862 134688 139890
rect 135272 139862 135516 139890
rect 136008 139862 136344 139890
rect 136744 139862 137172 139890
rect 137940 139862 138000 139890
rect 138584 139862 138828 139890
rect 139412 139862 139656 139890
rect 140148 139862 140484 139890
rect 140976 139862 141312 139890
rect 141436 139346 141464 177919
rect 141528 140185 141556 190426
rect 141712 148306 141740 190426
rect 142080 182034 142108 193186
rect 142160 193180 142212 193186
rect 142160 193122 142212 193128
rect 142264 191486 142292 198086
rect 142436 196444 142488 196450
rect 142436 196386 142488 196392
rect 142344 196104 142396 196110
rect 142344 196046 142396 196052
rect 142252 191480 142304 191486
rect 142252 191422 142304 191428
rect 142356 187338 142384 196046
rect 142448 192710 142476 196386
rect 142540 195022 142568 199650
rect 142632 197674 142660 199718
rect 142712 199708 142764 199714
rect 142712 199650 142764 199656
rect 142724 199510 142752 199650
rect 142712 199504 142764 199510
rect 142712 199446 142764 199452
rect 142908 199288 142936 199718
rect 142816 199260 142936 199288
rect 142712 198892 142764 198898
rect 142712 198834 142764 198840
rect 142724 198801 142752 198834
rect 142710 198792 142766 198801
rect 142710 198727 142766 198736
rect 142620 197668 142672 197674
rect 142620 197610 142672 197616
rect 142816 196110 142844 199260
rect 143000 199186 143028 199736
rect 143080 199640 143132 199646
rect 143080 199582 143132 199588
rect 142908 199158 143028 199186
rect 142804 196104 142856 196110
rect 142804 196046 142856 196052
rect 142908 195974 142936 199158
rect 142988 199096 143040 199102
rect 143092 199073 143120 199582
rect 142988 199038 143040 199044
rect 143078 199064 143134 199073
rect 143000 198801 143028 199038
rect 143078 198999 143134 199008
rect 142986 198792 143042 198801
rect 142986 198727 143042 198736
rect 143080 198552 143132 198558
rect 143080 198494 143132 198500
rect 142632 195946 142936 195974
rect 142528 195016 142580 195022
rect 142528 194958 142580 194964
rect 142528 194880 142580 194886
rect 142528 194822 142580 194828
rect 142436 192704 142488 192710
rect 142436 192646 142488 192652
rect 142344 187332 142396 187338
rect 142344 187274 142396 187280
rect 142068 182028 142120 182034
rect 142068 181970 142120 181976
rect 142448 181558 142476 192646
rect 142436 181552 142488 181558
rect 142436 181494 142488 181500
rect 142540 180577 142568 194822
rect 142526 180568 142582 180577
rect 142526 180503 142582 180512
rect 142540 180033 142568 180503
rect 142526 180024 142582 180033
rect 142526 179959 142582 179968
rect 142632 148578 142660 195946
rect 143092 195242 143120 198494
rect 143184 196722 143212 199736
rect 143262 199744 143350 199753
rect 143318 199736 143350 199744
rect 143414 199764 143442 200124
rect 143506 199918 143534 200124
rect 143494 199912 143546 199918
rect 143494 199854 143546 199860
rect 143598 199764 143626 200124
rect 143414 199736 143488 199764
rect 143262 199679 143318 199688
rect 143460 199617 143488 199736
rect 143552 199736 143626 199764
rect 143446 199608 143502 199617
rect 143446 199543 143502 199552
rect 143448 199504 143500 199510
rect 143448 199446 143500 199452
rect 143460 198150 143488 199446
rect 143448 198144 143500 198150
rect 143448 198086 143500 198092
rect 143448 198008 143500 198014
rect 143448 197950 143500 197956
rect 143354 196752 143410 196761
rect 143172 196716 143224 196722
rect 143354 196687 143410 196696
rect 143172 196658 143224 196664
rect 143170 195936 143226 195945
rect 143170 195871 143226 195880
rect 142816 195214 143120 195242
rect 142816 189650 142844 195214
rect 142986 195120 143042 195129
rect 142986 195055 143042 195064
rect 143000 193118 143028 195055
rect 142988 193112 143040 193118
rect 142988 193054 143040 193060
rect 143184 191834 143212 195871
rect 143000 191806 143212 191834
rect 142804 189644 142856 189650
rect 142804 189586 142856 189592
rect 142804 188012 142856 188018
rect 142804 187954 142856 187960
rect 142620 148572 142672 148578
rect 142620 148514 142672 148520
rect 142816 148481 142844 187954
rect 143000 187105 143028 191806
rect 143368 187202 143396 196687
rect 143460 188970 143488 197950
rect 143552 196790 143580 199736
rect 143690 199696 143718 200124
rect 143782 199918 143810 200124
rect 143770 199912 143822 199918
rect 143770 199854 143822 199860
rect 143874 199764 143902 200124
rect 143644 199668 143718 199696
rect 143828 199736 143902 199764
rect 143540 196784 143592 196790
rect 143540 196726 143592 196732
rect 143644 196602 143672 199668
rect 143724 199572 143776 199578
rect 143724 199514 143776 199520
rect 143736 196722 143764 199514
rect 143828 197402 143856 199736
rect 143966 199696 143994 200124
rect 144058 199918 144086 200124
rect 144046 199912 144098 199918
rect 144046 199854 144098 199860
rect 143920 199668 143994 199696
rect 144150 199696 144178 200124
rect 144242 199764 144270 200124
rect 144334 199918 144362 200124
rect 144322 199912 144374 199918
rect 144322 199854 144374 199860
rect 144426 199764 144454 200124
rect 144518 199889 144546 200124
rect 144504 199880 144560 199889
rect 144504 199815 144560 199824
rect 144610 199764 144638 200124
rect 144702 199918 144730 200124
rect 144794 199918 144822 200124
rect 144690 199912 144742 199918
rect 144690 199854 144742 199860
rect 144782 199912 144834 199918
rect 144782 199854 144834 199860
rect 144886 199764 144914 200124
rect 144242 199736 144316 199764
rect 144150 199668 144224 199696
rect 143816 197396 143868 197402
rect 143816 197338 143868 197344
rect 143724 196716 143776 196722
rect 143724 196658 143776 196664
rect 143644 196574 143856 196602
rect 143724 196512 143776 196518
rect 143724 196454 143776 196460
rect 143448 188964 143500 188970
rect 143448 188906 143500 188912
rect 143448 188828 143500 188834
rect 143448 188770 143500 188776
rect 143460 188737 143488 188770
rect 143446 188728 143502 188737
rect 143446 188663 143502 188672
rect 143460 187814 143488 188663
rect 143448 187808 143500 187814
rect 143448 187750 143500 187756
rect 143356 187196 143408 187202
rect 143356 187138 143408 187144
rect 142986 187096 143042 187105
rect 142986 187031 143042 187040
rect 143736 184278 143764 196454
rect 143828 184890 143856 196574
rect 143816 184884 143868 184890
rect 143816 184826 143868 184832
rect 143920 184346 143948 199668
rect 144000 199572 144052 199578
rect 144000 199514 144052 199520
rect 144012 198694 144040 199514
rect 144092 199504 144144 199510
rect 144092 199446 144144 199452
rect 144104 199209 144132 199446
rect 144090 199200 144146 199209
rect 144090 199135 144146 199144
rect 144000 198688 144052 198694
rect 144000 198630 144052 198636
rect 144196 198472 144224 199668
rect 144012 198444 144224 198472
rect 144012 195537 144040 198444
rect 144092 198348 144144 198354
rect 144092 198290 144144 198296
rect 143998 195528 144054 195537
rect 143998 195463 144054 195472
rect 144000 195424 144052 195430
rect 144000 195366 144052 195372
rect 143908 184340 143960 184346
rect 143908 184282 143960 184288
rect 143724 184272 143776 184278
rect 143724 184214 143776 184220
rect 143446 182200 143502 182209
rect 143446 182135 143448 182144
rect 143500 182135 143502 182144
rect 143448 182106 143500 182112
rect 142802 148472 142858 148481
rect 144012 148442 144040 195366
rect 144104 192370 144132 198290
rect 144184 197940 144236 197946
rect 144184 197882 144236 197888
rect 144196 195430 144224 197882
rect 144288 196874 144316 199736
rect 144380 199736 144454 199764
rect 144564 199736 144638 199764
rect 144840 199736 144914 199764
rect 144380 197169 144408 199736
rect 144460 199640 144512 199646
rect 144460 199582 144512 199588
rect 144472 197606 144500 199582
rect 144564 198762 144592 199736
rect 144736 199708 144788 199714
rect 144736 199650 144788 199656
rect 144748 199617 144776 199650
rect 144734 199608 144790 199617
rect 144644 199572 144696 199578
rect 144734 199543 144790 199552
rect 144644 199514 144696 199520
rect 144552 198756 144604 198762
rect 144552 198698 144604 198704
rect 144460 197600 144512 197606
rect 144460 197542 144512 197548
rect 144366 197160 144422 197169
rect 144366 197095 144422 197104
rect 144288 196846 144592 196874
rect 144460 196784 144512 196790
rect 144460 196726 144512 196732
rect 144276 196716 144328 196722
rect 144276 196658 144328 196664
rect 144184 195424 144236 195430
rect 144184 195366 144236 195372
rect 144182 194576 144238 194585
rect 144182 194511 144238 194520
rect 144092 192364 144144 192370
rect 144092 192306 144144 192312
rect 144196 186386 144224 194511
rect 144288 191826 144316 196658
rect 144276 191820 144328 191826
rect 144276 191762 144328 191768
rect 144184 186380 144236 186386
rect 144184 186322 144236 186328
rect 144182 183424 144238 183433
rect 144182 183359 144238 183368
rect 144196 182753 144224 183359
rect 144182 182744 144238 182753
rect 144182 182679 144238 182688
rect 142802 148407 142858 148416
rect 144000 148436 144052 148442
rect 144000 148378 144052 148384
rect 141700 148300 141752 148306
rect 141700 148242 141752 148248
rect 144092 145852 144144 145858
rect 144092 145794 144144 145800
rect 141792 144696 141844 144702
rect 141792 144638 141844 144644
rect 141514 140176 141570 140185
rect 141514 140111 141570 140120
rect 141804 139890 141832 144638
rect 142896 144628 142948 144634
rect 142896 144570 142948 144576
rect 142908 142458 142936 144570
rect 143540 143064 143592 143070
rect 143540 143006 143592 143012
rect 142896 142452 142948 142458
rect 142896 142394 142948 142400
rect 142908 139890 142936 142394
rect 143552 139890 143580 143006
rect 144104 142154 144132 145794
rect 144196 144401 144224 182679
rect 144472 148782 144500 196726
rect 144564 183938 144592 196846
rect 144656 196518 144684 199514
rect 144736 199504 144788 199510
rect 144736 199446 144788 199452
rect 144748 199073 144776 199446
rect 144734 199064 144790 199073
rect 144734 198999 144790 199008
rect 144840 198734 144868 199736
rect 144978 199696 145006 200124
rect 145070 199918 145098 200124
rect 145058 199912 145110 199918
rect 145058 199854 145110 199860
rect 144748 198706 144868 198734
rect 144932 199668 145006 199696
rect 144748 196586 144776 198706
rect 144828 196920 144880 196926
rect 144828 196862 144880 196868
rect 144736 196580 144788 196586
rect 144736 196522 144788 196528
rect 144644 196512 144696 196518
rect 144644 196454 144696 196460
rect 144840 192302 144868 196862
rect 144932 196450 144960 199668
rect 145162 199594 145190 200124
rect 145254 199850 145282 200124
rect 145242 199844 145294 199850
rect 145242 199786 145294 199792
rect 145346 199730 145374 200124
rect 145438 199918 145466 200124
rect 145530 199918 145558 200124
rect 145622 199918 145650 200124
rect 145426 199912 145478 199918
rect 145426 199854 145478 199860
rect 145518 199912 145570 199918
rect 145518 199854 145570 199860
rect 145610 199912 145662 199918
rect 145610 199854 145662 199860
rect 145714 199764 145742 200124
rect 145806 199889 145834 200124
rect 145898 199918 145926 200124
rect 145886 199912 145938 199918
rect 145792 199880 145848 199889
rect 145886 199854 145938 199860
rect 145792 199815 145848 199824
rect 145714 199736 145788 199764
rect 145012 199572 145064 199578
rect 145012 199514 145064 199520
rect 145116 199566 145190 199594
rect 145300 199702 145374 199730
rect 145472 199708 145524 199714
rect 144920 196444 144972 196450
rect 144920 196386 144972 196392
rect 145024 194585 145052 199514
rect 145116 198354 145144 199566
rect 145196 199096 145248 199102
rect 145196 199038 145248 199044
rect 145208 198898 145236 199038
rect 145196 198892 145248 198898
rect 145196 198834 145248 198840
rect 145104 198348 145156 198354
rect 145104 198290 145156 198296
rect 145300 196704 145328 199702
rect 145472 199650 145524 199656
rect 145564 199708 145616 199714
rect 145564 199650 145616 199656
rect 145380 199640 145432 199646
rect 145380 199582 145432 199588
rect 145116 196676 145328 196704
rect 145010 194576 145066 194585
rect 145010 194511 145066 194520
rect 144828 192296 144880 192302
rect 144828 192238 144880 192244
rect 144644 189032 144696 189038
rect 144642 189000 144644 189009
rect 144696 189000 144698 189009
rect 144642 188935 144698 188944
rect 144656 187746 144684 188935
rect 144644 187740 144696 187746
rect 144644 187682 144696 187688
rect 145116 187270 145144 196676
rect 145196 196580 145248 196586
rect 145196 196522 145248 196528
rect 145208 188358 145236 196522
rect 145392 195158 145420 199582
rect 145380 195152 145432 195158
rect 145380 195094 145432 195100
rect 145196 188352 145248 188358
rect 145196 188294 145248 188300
rect 145104 187264 145156 187270
rect 145104 187206 145156 187212
rect 144828 186380 144880 186386
rect 144828 186322 144880 186328
rect 144734 186280 144790 186289
rect 144734 186215 144790 186224
rect 144748 184890 144776 186215
rect 144840 186182 144868 186322
rect 144828 186176 144880 186182
rect 144828 186118 144880 186124
rect 144736 184884 144788 184890
rect 144736 184826 144788 184832
rect 144748 184210 144776 184826
rect 144828 184816 144880 184822
rect 144828 184758 144880 184764
rect 144840 184278 144868 184758
rect 144828 184272 144880 184278
rect 144828 184214 144880 184220
rect 144736 184204 144788 184210
rect 144736 184146 144788 184152
rect 144552 183932 144604 183938
rect 144552 183874 144604 183880
rect 144460 148776 144512 148782
rect 144460 148718 144512 148724
rect 144182 144392 144238 144401
rect 144182 144327 144238 144336
rect 145196 144356 145248 144362
rect 145196 144298 145248 144304
rect 144104 142126 144224 142154
rect 144196 139890 144224 142126
rect 145208 139890 145236 144298
rect 145484 140282 145512 199650
rect 145576 198734 145604 199650
rect 145656 199300 145708 199306
rect 145656 199242 145708 199248
rect 145668 198898 145696 199242
rect 145656 198892 145708 198898
rect 145656 198834 145708 198840
rect 145576 198706 145696 198734
rect 145564 197804 145616 197810
rect 145564 197746 145616 197752
rect 145576 141370 145604 197746
rect 145668 186318 145696 198706
rect 145760 193050 145788 199736
rect 145990 199730 146018 200124
rect 145944 199702 146018 199730
rect 145840 199368 145892 199374
rect 145840 199310 145892 199316
rect 145852 196586 145880 199310
rect 145944 197878 145972 199702
rect 146082 199594 146110 200124
rect 146174 199764 146202 200124
rect 146266 199918 146294 200124
rect 146358 199918 146386 200124
rect 146450 199923 146478 200124
rect 146254 199912 146306 199918
rect 146254 199854 146306 199860
rect 146346 199912 146398 199918
rect 146346 199854 146398 199860
rect 146436 199914 146492 199923
rect 146542 199918 146570 200124
rect 146436 199849 146492 199858
rect 146530 199912 146582 199918
rect 146530 199854 146582 199860
rect 146634 199850 146662 200124
rect 146726 199923 146754 200124
rect 146712 199914 146768 199923
rect 146818 199918 146846 200124
rect 146910 199918 146938 200124
rect 146622 199844 146674 199850
rect 146712 199849 146768 199858
rect 146806 199912 146858 199918
rect 146806 199854 146858 199860
rect 146898 199912 146950 199918
rect 146898 199854 146950 199860
rect 147002 199850 147030 200124
rect 147094 199923 147122 200124
rect 147080 199914 147136 199923
rect 147186 199918 147214 200124
rect 147278 199918 147306 200124
rect 147370 199923 147398 200124
rect 146622 199786 146674 199792
rect 146990 199844 147042 199850
rect 147080 199849 147136 199858
rect 147174 199912 147226 199918
rect 147174 199854 147226 199860
rect 147266 199912 147318 199918
rect 147266 199854 147318 199860
rect 147356 199914 147412 199923
rect 147356 199849 147412 199858
rect 146990 199786 147042 199792
rect 147462 199764 147490 200124
rect 146174 199736 146248 199764
rect 146036 199566 146110 199594
rect 146036 198558 146064 199566
rect 146024 198552 146076 198558
rect 146024 198494 146076 198500
rect 145932 197872 145984 197878
rect 145932 197814 145984 197820
rect 146220 197713 146248 199736
rect 146850 199744 146906 199753
rect 146484 199708 146536 199714
rect 146484 199650 146536 199656
rect 146668 199708 146720 199714
rect 147034 199744 147090 199753
rect 146850 199679 146906 199688
rect 146944 199708 146996 199714
rect 146668 199650 146720 199656
rect 146392 199640 146444 199646
rect 146392 199582 146444 199588
rect 146300 199572 146352 199578
rect 146300 199514 146352 199520
rect 146206 197704 146262 197713
rect 146206 197639 146262 197648
rect 146312 197282 146340 199514
rect 146220 197254 146340 197282
rect 146114 197160 146170 197169
rect 146114 197095 146170 197104
rect 146128 196625 146156 197095
rect 146114 196616 146170 196625
rect 145840 196580 145892 196586
rect 146114 196551 146170 196560
rect 145840 196522 145892 196528
rect 145840 196444 145892 196450
rect 145840 196386 145892 196392
rect 145748 193044 145800 193050
rect 145748 192986 145800 192992
rect 145852 190126 145880 196386
rect 146220 194070 146248 197254
rect 146404 196790 146432 199582
rect 146392 196784 146444 196790
rect 146392 196726 146444 196732
rect 146496 194594 146524 199650
rect 146574 199608 146630 199617
rect 146574 199543 146576 199552
rect 146628 199543 146630 199552
rect 146576 199514 146628 199520
rect 146576 199300 146628 199306
rect 146576 199242 146628 199248
rect 146312 194566 146524 194594
rect 146208 194064 146260 194070
rect 146208 194006 146260 194012
rect 146208 193928 146260 193934
rect 146208 193870 146260 193876
rect 145840 190120 145892 190126
rect 145840 190062 145892 190068
rect 145656 186312 145708 186318
rect 145656 186254 145708 186260
rect 146220 147914 146248 193870
rect 146312 192778 146340 194566
rect 146300 192772 146352 192778
rect 146300 192714 146352 192720
rect 146588 190194 146616 199242
rect 146680 197402 146708 199650
rect 146760 199640 146812 199646
rect 146760 199582 146812 199588
rect 146772 197470 146800 199582
rect 146760 197464 146812 197470
rect 146760 197406 146812 197412
rect 146668 197396 146720 197402
rect 146668 197338 146720 197344
rect 146668 197124 146720 197130
rect 146668 197066 146720 197072
rect 146680 193866 146708 197066
rect 146864 196874 146892 199679
rect 147034 199679 147090 199688
rect 147416 199736 147490 199764
rect 147554 199764 147582 200124
rect 147646 199918 147674 200124
rect 147738 199918 147766 200124
rect 147634 199912 147686 199918
rect 147634 199854 147686 199860
rect 147726 199912 147778 199918
rect 147726 199854 147778 199860
rect 147830 199764 147858 200124
rect 147922 199918 147950 200124
rect 148014 199918 148042 200124
rect 148106 199918 148134 200124
rect 148198 199923 148226 200124
rect 147910 199912 147962 199918
rect 147910 199854 147962 199860
rect 148002 199912 148054 199918
rect 148002 199854 148054 199860
rect 148094 199912 148146 199918
rect 148094 199854 148146 199860
rect 148184 199914 148240 199923
rect 148290 199918 148318 200124
rect 148184 199849 148240 199858
rect 148278 199912 148330 199918
rect 148278 199854 148330 199860
rect 147554 199736 147628 199764
rect 146944 199650 146996 199656
rect 146956 198014 146984 199650
rect 146944 198008 146996 198014
rect 146944 197950 146996 197956
rect 147048 196926 147076 199679
rect 147220 199640 147272 199646
rect 147220 199582 147272 199588
rect 147310 199608 147366 199617
rect 147128 197396 147180 197402
rect 147128 197338 147180 197344
rect 147036 196920 147088 196926
rect 146864 196846 146984 196874
rect 147036 196862 147088 196868
rect 146852 196784 146904 196790
rect 146956 196772 146984 196846
rect 146956 196744 147076 196772
rect 146852 196726 146904 196732
rect 146760 196716 146812 196722
rect 146760 196658 146812 196664
rect 146668 193860 146720 193866
rect 146668 193802 146720 193808
rect 146666 193760 146722 193769
rect 146666 193695 146722 193704
rect 146576 190188 146628 190194
rect 146576 190130 146628 190136
rect 146220 147886 146340 147914
rect 146312 147801 146340 147886
rect 146298 147792 146354 147801
rect 146298 147727 146354 147736
rect 146312 144294 146340 147727
rect 146300 144288 146352 144294
rect 146300 144230 146352 144236
rect 145932 143132 145984 143138
rect 145932 143074 145984 143080
rect 145564 141364 145616 141370
rect 145564 141306 145616 141312
rect 145472 140276 145524 140282
rect 145472 140218 145524 140224
rect 145944 139890 145972 143074
rect 146680 142050 146708 193695
rect 146772 187134 146800 196658
rect 146864 190262 146892 196726
rect 146942 196616 146998 196625
rect 146942 196551 146998 196560
rect 146852 190256 146904 190262
rect 146852 190198 146904 190204
rect 146760 187128 146812 187134
rect 146760 187070 146812 187076
rect 146758 142760 146814 142769
rect 146758 142695 146814 142704
rect 146668 142044 146720 142050
rect 146668 141986 146720 141992
rect 146668 140004 146720 140010
rect 146668 139946 146720 139952
rect 141804 139862 142140 139890
rect 142908 139862 142968 139890
rect 143552 139862 143796 139890
rect 144196 139862 144624 139890
rect 145208 139862 145452 139890
rect 145944 139862 146280 139890
rect 146680 139369 146708 139946
rect 146772 139890 146800 142695
rect 146956 140010 146984 196551
rect 147048 187406 147076 196744
rect 147140 194313 147168 197338
rect 147232 195702 147260 199582
rect 147310 199543 147366 199552
rect 147324 198529 147352 199543
rect 147310 198520 147366 198529
rect 147310 198455 147366 198464
rect 147416 198393 147444 199736
rect 147496 199640 147548 199646
rect 147496 199582 147548 199588
rect 147402 198384 147458 198393
rect 147402 198319 147458 198328
rect 147312 197464 147364 197470
rect 147312 197406 147364 197412
rect 147220 195696 147272 195702
rect 147220 195638 147272 195644
rect 147126 194304 147182 194313
rect 147126 194239 147182 194248
rect 147140 192386 147168 194239
rect 147324 193214 147352 197406
rect 147232 193186 147352 193214
rect 147232 192506 147260 193186
rect 147508 192817 147536 199582
rect 147600 196722 147628 199736
rect 147784 199736 147858 199764
rect 147956 199776 148008 199782
rect 147680 199708 147732 199714
rect 147680 199650 147732 199656
rect 147692 196722 147720 199650
rect 147588 196716 147640 196722
rect 147588 196658 147640 196664
rect 147680 196716 147732 196722
rect 147680 196658 147732 196664
rect 147784 195702 147812 199736
rect 147956 199718 148008 199724
rect 147864 199640 147916 199646
rect 147862 199608 147864 199617
rect 147916 199608 147918 199617
rect 147862 199543 147918 199552
rect 147864 199504 147916 199510
rect 147864 199446 147916 199452
rect 147876 197538 147904 199446
rect 147968 199034 147996 199718
rect 148232 199708 148284 199714
rect 148232 199650 148284 199656
rect 148140 199640 148192 199646
rect 148140 199582 148192 199588
rect 148048 199572 148100 199578
rect 148048 199514 148100 199520
rect 147956 199028 148008 199034
rect 147956 198970 148008 198976
rect 147956 198416 148008 198422
rect 147956 198358 148008 198364
rect 147968 198132 147996 198358
rect 148060 198286 148088 199514
rect 148048 198280 148100 198286
rect 148048 198222 148100 198228
rect 147968 198104 148088 198132
rect 148060 197674 148088 198104
rect 148048 197668 148100 197674
rect 148048 197610 148100 197616
rect 147864 197532 147916 197538
rect 147864 197474 147916 197480
rect 147956 197396 148008 197402
rect 147956 197338 148008 197344
rect 147772 195696 147824 195702
rect 147772 195638 147824 195644
rect 147680 193452 147732 193458
rect 147680 193394 147732 193400
rect 147586 192944 147642 192953
rect 147586 192879 147642 192888
rect 147494 192808 147550 192817
rect 147494 192743 147550 192752
rect 147220 192500 147272 192506
rect 147220 192442 147272 192448
rect 147140 192358 147260 192386
rect 147036 187400 147088 187406
rect 147036 187342 147088 187348
rect 147232 187241 147260 192358
rect 147310 189136 147366 189145
rect 147310 189071 147366 189080
rect 147218 187232 147274 187241
rect 147218 187167 147274 187176
rect 147324 140049 147352 189071
rect 147600 185638 147628 192879
rect 147692 192846 147720 193394
rect 147680 192840 147732 192846
rect 147680 192782 147732 192788
rect 147588 185632 147640 185638
rect 147588 185574 147640 185580
rect 147968 180794 147996 197338
rect 148060 190454 148088 197610
rect 148152 197130 148180 199582
rect 148244 197810 148272 199650
rect 148382 199458 148410 200124
rect 148474 199850 148502 200124
rect 148566 199918 148594 200124
rect 148658 199918 148686 200124
rect 148554 199912 148606 199918
rect 148554 199854 148606 199860
rect 148646 199912 148698 199918
rect 148646 199854 148698 199860
rect 148462 199844 148514 199850
rect 148462 199786 148514 199792
rect 148750 199753 148778 200124
rect 148842 199782 148870 200124
rect 148934 199918 148962 200124
rect 148922 199912 148974 199918
rect 149026 199889 149054 200124
rect 149118 199918 149146 200124
rect 149106 199912 149158 199918
rect 148922 199854 148974 199860
rect 149012 199880 149068 199889
rect 149106 199854 149158 199860
rect 149012 199815 149068 199824
rect 148830 199776 148882 199782
rect 148736 199744 148792 199753
rect 148830 199718 148882 199724
rect 148968 199776 149020 199782
rect 148968 199718 149020 199724
rect 149058 199744 149114 199753
rect 148736 199679 148792 199688
rect 148784 199572 148836 199578
rect 148784 199514 148836 199520
rect 148336 199430 148410 199458
rect 148232 197804 148284 197810
rect 148232 197746 148284 197752
rect 148140 197124 148192 197130
rect 148140 197066 148192 197072
rect 148336 196926 148364 199430
rect 148416 198280 148468 198286
rect 148416 198222 148468 198228
rect 148324 196920 148376 196926
rect 148324 196862 148376 196868
rect 148140 196784 148192 196790
rect 148140 196726 148192 196732
rect 148152 191049 148180 196726
rect 148230 196480 148286 196489
rect 148230 196415 148286 196424
rect 148244 195634 148272 196415
rect 148324 196036 148376 196042
rect 148324 195978 148376 195984
rect 148232 195628 148284 195634
rect 148232 195570 148284 195576
rect 148138 191040 148194 191049
rect 148138 190975 148194 190984
rect 148060 190426 148180 190454
rect 147876 180766 147996 180794
rect 147680 143268 147732 143274
rect 147680 143210 147732 143216
rect 147310 140040 147366 140049
rect 146944 140004 146996 140010
rect 147310 139975 147366 139984
rect 146944 139946 146996 139952
rect 147692 139890 147720 143210
rect 147876 140758 147904 180766
rect 148152 148345 148180 190426
rect 148138 148336 148194 148345
rect 148138 148271 148194 148280
rect 148336 141642 148364 195978
rect 148428 144498 148456 198222
rect 148690 197976 148746 197985
rect 148690 197911 148746 197920
rect 148508 196920 148560 196926
rect 148508 196862 148560 196868
rect 148520 195974 148548 196862
rect 148520 195946 148640 195974
rect 148508 195696 148560 195702
rect 148508 195638 148560 195644
rect 148520 193594 148548 195638
rect 148508 193588 148560 193594
rect 148508 193530 148560 193536
rect 148416 144492 148468 144498
rect 148416 144434 148468 144440
rect 148414 142896 148470 142905
rect 148414 142831 148470 142840
rect 148324 141636 148376 141642
rect 148324 141578 148376 141584
rect 147864 140752 147916 140758
rect 147864 140694 147916 140700
rect 148428 139890 148456 142831
rect 148520 141846 148548 193530
rect 148612 190454 148640 195946
rect 148704 192846 148732 197911
rect 148796 196790 148824 199514
rect 148876 199368 148928 199374
rect 148876 199310 148928 199316
rect 148888 197860 148916 199310
rect 148980 197985 149008 199718
rect 149058 199679 149114 199688
rect 149210 199696 149238 200124
rect 149302 199764 149330 200124
rect 149394 199918 149422 200124
rect 149382 199912 149434 199918
rect 149486 199889 149514 200124
rect 149382 199854 149434 199860
rect 149472 199880 149528 199889
rect 149472 199815 149528 199824
rect 149428 199776 149480 199782
rect 149302 199736 149376 199764
rect 148966 197976 149022 197985
rect 148966 197911 149022 197920
rect 148888 197832 149008 197860
rect 148784 196784 148836 196790
rect 148784 196726 148836 196732
rect 148876 196716 148928 196722
rect 148876 196658 148928 196664
rect 148692 192840 148744 192846
rect 148692 192782 148744 192788
rect 148612 190426 148824 190454
rect 148796 171834 148824 190426
rect 148784 171828 148836 171834
rect 148784 171770 148836 171776
rect 148888 144430 148916 196658
rect 148980 196042 149008 197832
rect 149072 197810 149100 199679
rect 149210 199668 149284 199696
rect 149256 199560 149284 199668
rect 149164 199532 149284 199560
rect 149060 197804 149112 197810
rect 149060 197746 149112 197752
rect 149060 197464 149112 197470
rect 149060 197406 149112 197412
rect 148968 196036 149020 196042
rect 148968 195978 149020 195984
rect 149072 191078 149100 197406
rect 149164 196761 149192 199532
rect 149244 197124 149296 197130
rect 149244 197066 149296 197072
rect 149150 196752 149206 196761
rect 149150 196687 149206 196696
rect 149256 195412 149284 197066
rect 149348 195566 149376 199736
rect 149578 199764 149606 200124
rect 149428 199718 149480 199724
rect 149532 199736 149606 199764
rect 149440 196874 149468 199718
rect 149532 196994 149560 199736
rect 149670 199696 149698 200124
rect 149624 199668 149698 199696
rect 149520 196988 149572 196994
rect 149624 196976 149652 199668
rect 149762 199628 149790 200124
rect 149854 199918 149882 200124
rect 149842 199912 149894 199918
rect 149842 199854 149894 199860
rect 149946 199730 149974 200124
rect 150038 199918 150066 200124
rect 150130 199918 150158 200124
rect 150222 199918 150250 200124
rect 150026 199912 150078 199918
rect 150026 199854 150078 199860
rect 150118 199912 150170 199918
rect 150118 199854 150170 199860
rect 150210 199912 150262 199918
rect 150314 199889 150342 200124
rect 150406 199918 150434 200124
rect 150394 199912 150446 199918
rect 150210 199854 150262 199860
rect 150300 199880 150356 199889
rect 150394 199854 150446 199860
rect 150300 199815 150356 199824
rect 149716 199600 149790 199628
rect 149900 199702 149974 199730
rect 150072 199776 150124 199782
rect 150072 199718 150124 199724
rect 150348 199776 150400 199782
rect 150348 199718 150400 199724
rect 149716 197130 149744 199600
rect 149796 199504 149848 199510
rect 149796 199446 149848 199452
rect 149808 197130 149836 199446
rect 149704 197124 149756 197130
rect 149704 197066 149756 197072
rect 149796 197124 149848 197130
rect 149796 197066 149848 197072
rect 149624 196948 149836 196976
rect 149520 196930 149572 196936
rect 149440 196846 149744 196874
rect 149520 196716 149572 196722
rect 149520 196658 149572 196664
rect 149336 195560 149388 195566
rect 149336 195502 149388 195508
rect 149256 195384 149468 195412
rect 149336 193996 149388 194002
rect 149336 193938 149388 193944
rect 149060 191072 149112 191078
rect 149060 191014 149112 191020
rect 149348 180266 149376 193938
rect 149440 181558 149468 195384
rect 149532 189718 149560 196658
rect 149612 195968 149664 195974
rect 149612 195910 149664 195916
rect 149520 189712 149572 189718
rect 149520 189654 149572 189660
rect 149520 188352 149572 188358
rect 149520 188294 149572 188300
rect 149428 181552 149480 181558
rect 149428 181494 149480 181500
rect 149336 180260 149388 180266
rect 149336 180202 149388 180208
rect 148876 144424 148928 144430
rect 148876 144366 148928 144372
rect 149532 144129 149560 188294
rect 149518 144120 149574 144129
rect 149518 144055 149574 144064
rect 149244 142928 149296 142934
rect 149244 142870 149296 142876
rect 148508 141840 148560 141846
rect 148508 141782 148560 141788
rect 149256 139890 149284 142870
rect 149624 140214 149652 195910
rect 149716 188902 149744 196846
rect 149704 188896 149756 188902
rect 149704 188838 149756 188844
rect 149716 188766 149744 188838
rect 149704 188760 149756 188766
rect 149704 188702 149756 188708
rect 149702 182064 149758 182073
rect 149702 181999 149758 182008
rect 149716 144265 149744 181999
rect 149702 144256 149758 144265
rect 149702 144191 149758 144200
rect 149808 141710 149836 196948
rect 149900 195974 149928 199702
rect 149980 199640 150032 199646
rect 149980 199582 150032 199588
rect 149888 195968 149940 195974
rect 149888 195910 149940 195916
rect 149992 194002 150020 199582
rect 150084 196722 150112 199718
rect 150164 199708 150216 199714
rect 150164 199650 150216 199656
rect 150072 196716 150124 196722
rect 150072 196658 150124 196664
rect 149980 193996 150032 194002
rect 149980 193938 150032 193944
rect 150176 180794 150204 199650
rect 150254 199608 150310 199617
rect 150254 199543 150256 199552
rect 150308 199543 150310 199552
rect 150256 199514 150308 199520
rect 150256 199232 150308 199238
rect 150254 199200 150256 199209
rect 150308 199200 150310 199209
rect 150254 199135 150310 199144
rect 150256 199096 150308 199102
rect 150256 199038 150308 199044
rect 150268 198694 150296 199038
rect 150256 198688 150308 198694
rect 150256 198630 150308 198636
rect 150360 197470 150388 199718
rect 150498 199594 150526 200124
rect 150590 199918 150618 200124
rect 150682 199923 150710 200124
rect 150578 199912 150630 199918
rect 150578 199854 150630 199860
rect 150668 199914 150724 199923
rect 150668 199849 150724 199858
rect 150774 199850 150802 200124
rect 150866 199918 150894 200124
rect 150854 199912 150906 199918
rect 150854 199854 150906 199860
rect 150762 199844 150814 199850
rect 150762 199786 150814 199792
rect 150624 199776 150676 199782
rect 150624 199718 150676 199724
rect 150498 199566 150572 199594
rect 150440 199232 150492 199238
rect 150440 199174 150492 199180
rect 150348 197464 150400 197470
rect 150348 197406 150400 197412
rect 150348 197124 150400 197130
rect 150348 197066 150400 197072
rect 150360 191282 150388 197066
rect 150452 191593 150480 199174
rect 150544 197441 150572 199566
rect 150530 197432 150586 197441
rect 150530 197367 150586 197376
rect 150532 196716 150584 196722
rect 150532 196658 150584 196664
rect 150438 191584 150494 191593
rect 150438 191519 150494 191528
rect 150348 191276 150400 191282
rect 150348 191218 150400 191224
rect 150544 189922 150572 196658
rect 150532 189916 150584 189922
rect 150532 189858 150584 189864
rect 150636 182170 150664 199718
rect 150958 199696 150986 200124
rect 150912 199668 150986 199696
rect 150714 199608 150770 199617
rect 150714 199543 150716 199552
rect 150768 199543 150770 199552
rect 150716 199514 150768 199520
rect 150808 199300 150860 199306
rect 150808 199242 150860 199248
rect 150714 199064 150770 199073
rect 150714 198999 150770 199008
rect 150728 198626 150756 198999
rect 150716 198620 150768 198626
rect 150716 198562 150768 198568
rect 150728 197402 150756 198562
rect 150820 197674 150848 199242
rect 150912 198734 150940 199668
rect 151050 199628 151078 200124
rect 151142 199782 151170 200124
rect 151130 199776 151182 199782
rect 151130 199718 151182 199724
rect 151234 199730 151262 200124
rect 151326 199918 151354 200124
rect 151418 199918 151446 200124
rect 151314 199912 151366 199918
rect 151314 199854 151366 199860
rect 151406 199912 151458 199918
rect 151406 199854 151458 199860
rect 151360 199776 151412 199782
rect 151234 199702 151308 199730
rect 151510 199753 151538 200124
rect 151602 199918 151630 200124
rect 151590 199912 151642 199918
rect 151590 199854 151642 199860
rect 151694 199850 151722 200124
rect 151682 199844 151734 199850
rect 151682 199786 151734 199792
rect 151360 199718 151412 199724
rect 151496 199744 151552 199753
rect 151050 199600 151124 199628
rect 150992 199504 151044 199510
rect 150992 199446 151044 199452
rect 151004 199073 151032 199446
rect 150990 199064 151046 199073
rect 150990 198999 151046 199008
rect 150912 198706 151032 198734
rect 151004 198529 151032 198706
rect 150990 198520 151046 198529
rect 150990 198455 151046 198464
rect 151096 198121 151124 199600
rect 151280 199510 151308 199702
rect 151176 199504 151228 199510
rect 151176 199446 151228 199452
rect 151268 199504 151320 199510
rect 151268 199446 151320 199452
rect 151082 198112 151138 198121
rect 151082 198047 151138 198056
rect 150808 197668 150860 197674
rect 150808 197610 150860 197616
rect 150716 197396 150768 197402
rect 150716 197338 150768 197344
rect 151082 196752 151138 196761
rect 151082 196687 151138 196696
rect 150716 196512 150768 196518
rect 150716 196454 150768 196460
rect 150728 185706 150756 196454
rect 150992 195152 151044 195158
rect 150992 195094 151044 195100
rect 151004 189854 151032 195094
rect 150992 189848 151044 189854
rect 150992 189790 151044 189796
rect 150898 189136 150954 189145
rect 150898 189071 150954 189080
rect 150912 188766 150940 189071
rect 150900 188760 150952 188766
rect 150900 188702 150952 188708
rect 150912 188018 150940 188702
rect 150900 188012 150952 188018
rect 150900 187954 150952 187960
rect 151096 187474 151124 196687
rect 151084 187468 151136 187474
rect 151084 187410 151136 187416
rect 151188 187377 151216 199446
rect 151372 196518 151400 199718
rect 151496 199679 151552 199688
rect 151636 199708 151688 199714
rect 151636 199650 151688 199656
rect 151648 199617 151676 199650
rect 151786 199628 151814 200124
rect 151878 199764 151906 200124
rect 151970 199923 151998 200124
rect 151956 199914 152012 199923
rect 151956 199849 152012 199858
rect 152062 199850 152090 200124
rect 152154 199923 152182 200124
rect 152140 199914 152196 199923
rect 152050 199844 152102 199850
rect 152140 199849 152196 199858
rect 152246 199850 152274 200124
rect 152338 199923 152366 200124
rect 152324 199914 152380 199923
rect 152430 199918 152458 200124
rect 152050 199786 152102 199792
rect 152234 199844 152286 199850
rect 152324 199849 152380 199858
rect 152418 199912 152470 199918
rect 152418 199854 152470 199860
rect 152234 199786 152286 199792
rect 152522 199764 152550 200124
rect 152614 199850 152642 200124
rect 152706 199889 152734 200124
rect 152692 199880 152748 199889
rect 152602 199844 152654 199850
rect 152798 199850 152826 200124
rect 152692 199815 152748 199824
rect 152786 199844 152838 199850
rect 152602 199786 152654 199792
rect 152786 199786 152838 199792
rect 151878 199753 151952 199764
rect 151878 199744 151966 199753
rect 151878 199736 151910 199744
rect 151910 199679 151966 199688
rect 152094 199744 152150 199753
rect 152370 199744 152426 199753
rect 152150 199702 152228 199730
rect 152094 199679 152150 199688
rect 152096 199640 152148 199646
rect 151450 199608 151506 199617
rect 151634 199608 151690 199617
rect 151450 199543 151506 199552
rect 151544 199572 151596 199578
rect 151464 196722 151492 199543
rect 151786 199600 151952 199628
rect 151634 199543 151690 199552
rect 151544 199514 151596 199520
rect 151452 196716 151504 196722
rect 151452 196658 151504 196664
rect 151360 196512 151412 196518
rect 151360 196454 151412 196460
rect 151556 193214 151584 199514
rect 151728 199504 151780 199510
rect 151728 199446 151780 199452
rect 151636 199368 151688 199374
rect 151636 199310 151688 199316
rect 151648 199073 151676 199310
rect 151634 199064 151690 199073
rect 151634 198999 151690 199008
rect 151634 198928 151690 198937
rect 151634 198863 151690 198872
rect 151648 198762 151676 198863
rect 151636 198756 151688 198762
rect 151636 198698 151688 198704
rect 151740 197713 151768 199446
rect 151924 199170 151952 199600
rect 152096 199582 152148 199588
rect 151912 199164 151964 199170
rect 151912 199106 151964 199112
rect 152108 199073 152136 199582
rect 152094 199064 152150 199073
rect 152094 198999 152150 199008
rect 151818 198928 151874 198937
rect 151818 198863 151874 198872
rect 151726 197704 151782 197713
rect 151726 197639 151782 197648
rect 151636 197532 151688 197538
rect 151636 197474 151688 197480
rect 151464 193186 151584 193214
rect 151174 187368 151230 187377
rect 151174 187303 151230 187312
rect 150716 185700 150768 185706
rect 150716 185642 150768 185648
rect 150624 182164 150676 182170
rect 150624 182106 150676 182112
rect 149900 180766 150204 180794
rect 149900 144566 149928 180766
rect 150070 145616 150126 145625
rect 150070 145551 150126 145560
rect 149888 144560 149940 144566
rect 149888 144502 149940 144508
rect 149796 141704 149848 141710
rect 149796 141646 149848 141652
rect 149612 140208 149664 140214
rect 149612 140150 149664 140156
rect 150084 139890 150112 145551
rect 150900 142996 150952 143002
rect 150900 142938 150952 142944
rect 150912 139890 150940 142938
rect 151464 142118 151492 193186
rect 151648 180794 151676 197474
rect 151832 193934 151860 198863
rect 152096 197872 152148 197878
rect 152096 197814 152148 197820
rect 152004 195492 152056 195498
rect 152004 195434 152056 195440
rect 151820 193928 151872 193934
rect 151820 193870 151872 193876
rect 152016 181626 152044 195434
rect 152108 190942 152136 197814
rect 152200 192778 152228 199702
rect 152476 199736 152550 199764
rect 152646 199744 152702 199753
rect 152476 199730 152504 199736
rect 152426 199702 152504 199730
rect 152370 199679 152426 199688
rect 152890 199730 152918 200124
rect 152982 199923 153010 200124
rect 152968 199914 153024 199923
rect 152968 199849 153024 199858
rect 153074 199764 153102 200124
rect 153166 199918 153194 200124
rect 153258 199918 153286 200124
rect 153154 199912 153206 199918
rect 153154 199854 153206 199860
rect 153246 199912 153298 199918
rect 153246 199854 153298 199860
rect 153350 199764 153378 200124
rect 153028 199736 153102 199764
rect 153258 199736 153378 199764
rect 152890 199714 152964 199730
rect 152890 199708 152976 199714
rect 152890 199702 152924 199708
rect 152646 199679 152702 199688
rect 152464 199640 152516 199646
rect 152464 199582 152516 199588
rect 152372 199504 152424 199510
rect 152372 199446 152424 199452
rect 152278 198928 152334 198937
rect 152278 198863 152334 198872
rect 152292 194041 152320 198863
rect 152278 194032 152334 194041
rect 152278 193967 152334 193976
rect 152188 192772 152240 192778
rect 152188 192714 152240 192720
rect 152096 190936 152148 190942
rect 152096 190878 152148 190884
rect 152004 181620 152056 181626
rect 152004 181562 152056 181568
rect 151556 180766 151676 180794
rect 151452 142112 151504 142118
rect 151452 142054 151504 142060
rect 151556 141982 151584 180766
rect 152384 151814 152412 199446
rect 152476 193662 152504 199582
rect 152660 199424 152688 199679
rect 152924 199650 152976 199656
rect 152832 199640 152884 199646
rect 152832 199582 152884 199588
rect 152922 199608 152978 199617
rect 152568 199396 152688 199424
rect 152464 193656 152516 193662
rect 152464 193598 152516 193604
rect 152476 189689 152504 193598
rect 152462 189680 152518 189689
rect 152462 189615 152518 189624
rect 152292 151786 152412 151814
rect 151912 145716 151964 145722
rect 151912 145658 151964 145664
rect 151544 141976 151596 141982
rect 151544 141918 151596 141924
rect 151924 140758 151952 145658
rect 152292 141778 152320 151786
rect 152568 148345 152596 199396
rect 152646 199200 152702 199209
rect 152646 199135 152702 199144
rect 152740 199164 152792 199170
rect 152660 199102 152688 199135
rect 152740 199106 152792 199112
rect 152648 199096 152700 199102
rect 152648 199038 152700 199044
rect 152752 198937 152780 199106
rect 152738 198928 152794 198937
rect 152738 198863 152794 198872
rect 152844 198336 152872 199582
rect 152922 199543 152978 199552
rect 152752 198308 152872 198336
rect 152646 196072 152702 196081
rect 152646 196007 152702 196016
rect 152660 194585 152688 196007
rect 152752 195158 152780 198308
rect 152936 198234 152964 199543
rect 152844 198206 152964 198234
rect 152844 196722 152872 198206
rect 152924 198144 152976 198150
rect 152924 198086 152976 198092
rect 152832 196716 152884 196722
rect 152832 196658 152884 196664
rect 152740 195152 152792 195158
rect 152740 195094 152792 195100
rect 152646 194576 152702 194585
rect 152646 194511 152702 194520
rect 152660 189825 152688 194511
rect 152740 192772 152792 192778
rect 152740 192714 152792 192720
rect 152646 189816 152702 189825
rect 152646 189751 152702 189760
rect 152752 188358 152780 192714
rect 152740 188352 152792 188358
rect 152740 188294 152792 188300
rect 152936 181830 152964 198086
rect 153028 195498 153056 199736
rect 153258 199560 153286 199736
rect 153442 199696 153470 200124
rect 153396 199668 153470 199696
rect 153534 199696 153562 200124
rect 153626 199923 153654 200124
rect 153612 199914 153668 199923
rect 153612 199849 153668 199858
rect 153718 199696 153746 200124
rect 153534 199668 153608 199696
rect 153396 199617 153424 199668
rect 153382 199608 153438 199617
rect 153258 199532 153332 199560
rect 153382 199543 153438 199552
rect 153476 199572 153528 199578
rect 153200 199436 153252 199442
rect 153200 199378 153252 199384
rect 153108 199232 153160 199238
rect 153106 199200 153108 199209
rect 153160 199200 153162 199209
rect 153106 199135 153162 199144
rect 153108 196988 153160 196994
rect 153108 196930 153160 196936
rect 153016 195492 153068 195498
rect 153016 195434 153068 195440
rect 153120 190398 153148 196930
rect 153212 194138 153240 199378
rect 153304 196489 153332 199532
rect 153476 199514 153528 199520
rect 153384 199436 153436 199442
rect 153384 199378 153436 199384
rect 153290 196480 153346 196489
rect 153290 196415 153346 196424
rect 153290 196208 153346 196217
rect 153396 196178 153424 199378
rect 153290 196143 153346 196152
rect 153384 196172 153436 196178
rect 153200 194132 153252 194138
rect 153200 194074 153252 194080
rect 153304 191214 153332 196143
rect 153384 196114 153436 196120
rect 153382 196072 153438 196081
rect 153382 196007 153438 196016
rect 153292 191208 153344 191214
rect 153292 191150 153344 191156
rect 153108 190392 153160 190398
rect 153108 190334 153160 190340
rect 153108 188556 153160 188562
rect 153108 188498 153160 188504
rect 153120 188426 153148 188498
rect 153108 188420 153160 188426
rect 153108 188362 153160 188368
rect 152924 181824 152976 181830
rect 152924 181766 152976 181772
rect 152554 148336 152610 148345
rect 152554 148271 152610 148280
rect 152372 145580 152424 145586
rect 152372 145522 152424 145528
rect 152384 142322 152412 145522
rect 152372 142316 152424 142322
rect 152372 142258 152424 142264
rect 152280 141772 152332 141778
rect 152280 141714 152332 141720
rect 151912 140752 151964 140758
rect 151912 140694 151964 140700
rect 152384 139890 152412 142258
rect 153120 141642 153148 188362
rect 153396 182850 153424 196007
rect 153488 186969 153516 199514
rect 153580 196194 153608 199668
rect 153672 199668 153746 199696
rect 153672 196296 153700 199668
rect 153810 199560 153838 200124
rect 153902 199918 153930 200124
rect 153994 199918 154022 200124
rect 154086 199918 154114 200124
rect 153890 199912 153942 199918
rect 153890 199854 153942 199860
rect 153982 199912 154034 199918
rect 153982 199854 154034 199860
rect 154074 199912 154126 199918
rect 154074 199854 154126 199860
rect 154028 199776 154080 199782
rect 153934 199744 153990 199753
rect 154178 199764 154206 200124
rect 154270 199918 154298 200124
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 154362 199764 154390 200124
rect 154454 199918 154482 200124
rect 154442 199912 154494 199918
rect 154546 199889 154574 200124
rect 154638 199918 154666 200124
rect 154730 199918 154758 200124
rect 154822 199918 154850 200124
rect 154914 199918 154942 200124
rect 155006 199918 155034 200124
rect 154626 199912 154678 199918
rect 154442 199854 154494 199860
rect 154532 199880 154588 199889
rect 154626 199854 154678 199860
rect 154718 199912 154770 199918
rect 154718 199854 154770 199860
rect 154810 199912 154862 199918
rect 154810 199854 154862 199860
rect 154902 199912 154954 199918
rect 154902 199854 154954 199860
rect 154994 199912 155046 199918
rect 154994 199854 155046 199860
rect 154532 199815 154588 199824
rect 155098 199764 155126 200124
rect 154028 199718 154080 199724
rect 154132 199736 154206 199764
rect 154316 199736 154390 199764
rect 155052 199736 155126 199764
rect 153934 199679 153990 199688
rect 153764 199532 153838 199560
rect 153764 199442 153792 199532
rect 153752 199436 153804 199442
rect 153752 199378 153804 199384
rect 153844 199436 153896 199442
rect 153844 199378 153896 199384
rect 153750 198928 153806 198937
rect 153750 198863 153806 198872
rect 153764 196432 153792 198863
rect 153856 196994 153884 199378
rect 153948 199209 153976 199679
rect 153934 199200 153990 199209
rect 154040 199170 154068 199718
rect 153934 199135 153990 199144
rect 154028 199164 154080 199170
rect 153948 197538 153976 199135
rect 154028 199106 154080 199112
rect 153936 197532 153988 197538
rect 153936 197474 153988 197480
rect 153844 196988 153896 196994
rect 153844 196930 153896 196936
rect 153764 196404 153884 196432
rect 153672 196268 153792 196296
rect 153580 196166 153700 196194
rect 153568 196104 153620 196110
rect 153568 196046 153620 196052
rect 153580 189009 153608 196046
rect 153672 189689 153700 196166
rect 153658 189680 153714 189689
rect 153658 189615 153714 189624
rect 153566 189000 153622 189009
rect 153566 188935 153622 188944
rect 153580 188601 153608 188935
rect 153566 188592 153622 188601
rect 153566 188527 153622 188536
rect 153474 186960 153530 186969
rect 153474 186895 153530 186904
rect 153384 182844 153436 182850
rect 153384 182786 153436 182792
rect 153764 145790 153792 196268
rect 153856 195537 153884 196404
rect 153842 195528 153898 195537
rect 153842 195463 153898 195472
rect 154132 193769 154160 199736
rect 154212 199640 154264 199646
rect 154212 199582 154264 199588
rect 154224 195702 154252 199582
rect 154212 195696 154264 195702
rect 154212 195638 154264 195644
rect 154118 193760 154174 193769
rect 154118 193695 154174 193704
rect 154316 180794 154344 199736
rect 154488 199708 154540 199714
rect 154488 199650 154540 199656
rect 154580 199708 154632 199714
rect 154580 199650 154632 199656
rect 154672 199708 154724 199714
rect 154672 199650 154724 199656
rect 154764 199708 154816 199714
rect 154764 199650 154816 199656
rect 154856 199708 154908 199714
rect 154856 199650 154908 199656
rect 154396 199640 154448 199646
rect 154394 199608 154396 199617
rect 154448 199608 154450 199617
rect 154394 199543 154450 199552
rect 154500 196081 154528 199650
rect 154592 196874 154620 199650
rect 154684 198150 154712 199650
rect 154672 198144 154724 198150
rect 154672 198086 154724 198092
rect 154776 197878 154804 199650
rect 154868 198694 154896 199650
rect 154948 199368 155000 199374
rect 154948 199310 155000 199316
rect 154960 199102 154988 199310
rect 154948 199096 155000 199102
rect 154948 199038 155000 199044
rect 154856 198688 154908 198694
rect 154856 198630 154908 198636
rect 154764 197872 154816 197878
rect 154764 197814 154816 197820
rect 154960 197538 154988 199038
rect 154948 197532 155000 197538
rect 154948 197474 155000 197480
rect 154592 196846 154804 196874
rect 154672 196784 154724 196790
rect 154672 196726 154724 196732
rect 154486 196072 154542 196081
rect 154486 196007 154542 196016
rect 154488 195696 154540 195702
rect 154488 195638 154540 195644
rect 154500 191350 154528 195638
rect 154488 191344 154540 191350
rect 154488 191286 154540 191292
rect 154396 188488 154448 188494
rect 154396 188430 154448 188436
rect 154408 187814 154436 188430
rect 154396 187808 154448 187814
rect 154396 187750 154448 187756
rect 153948 180766 154344 180794
rect 153948 151814 153976 180766
rect 153948 151786 154068 151814
rect 153752 145784 153804 145790
rect 153752 145726 153804 145732
rect 153384 142860 153436 142866
rect 153384 142802 153436 142808
rect 153108 141636 153160 141642
rect 153108 141578 153160 141584
rect 152556 140752 152608 140758
rect 152556 140694 152608 140700
rect 146772 139862 147108 139890
rect 147692 139862 147936 139890
rect 148428 139862 148764 139890
rect 149256 139862 149592 139890
rect 150084 139862 150420 139890
rect 150912 139862 151248 139890
rect 152076 139862 152412 139890
rect 152568 139890 152596 140694
rect 153396 139890 153424 142802
rect 152568 139862 152904 139890
rect 153396 139862 153732 139890
rect 154040 139369 154068 151786
rect 154408 140049 154436 187750
rect 154488 145648 154540 145654
rect 154488 145590 154540 145596
rect 154500 142594 154528 145590
rect 154488 142588 154540 142594
rect 154488 142530 154540 142536
rect 154394 140040 154450 140049
rect 154394 139975 154450 139984
rect 154500 139890 154528 142530
rect 154684 140146 154712 196726
rect 154776 151162 154804 196846
rect 154856 196580 154908 196586
rect 154856 196522 154908 196528
rect 154868 184482 154896 196522
rect 155052 196518 155080 199736
rect 155190 199696 155218 200124
rect 155282 199764 155310 200124
rect 155374 199918 155402 200124
rect 155362 199912 155414 199918
rect 155362 199854 155414 199860
rect 155466 199764 155494 200124
rect 155282 199736 155356 199764
rect 155144 199668 155218 199696
rect 155040 196512 155092 196518
rect 155040 196454 155092 196460
rect 155144 187814 155172 199668
rect 155224 199504 155276 199510
rect 155224 199446 155276 199452
rect 155236 198762 155264 199446
rect 155224 198756 155276 198762
rect 155224 198698 155276 198704
rect 155328 191418 155356 199736
rect 155420 199736 155494 199764
rect 155558 199764 155586 200124
rect 155650 199918 155678 200124
rect 155742 199918 155770 200124
rect 155834 199923 155862 200124
rect 155638 199912 155690 199918
rect 155638 199854 155690 199860
rect 155730 199912 155782 199918
rect 155730 199854 155782 199860
rect 155820 199914 155876 199923
rect 155820 199849 155876 199858
rect 155684 199776 155736 199782
rect 155558 199736 155632 199764
rect 155420 197656 155448 199736
rect 155500 199640 155552 199646
rect 155500 199582 155552 199588
rect 155512 199170 155540 199582
rect 155500 199164 155552 199170
rect 155500 199106 155552 199112
rect 155420 197628 155540 197656
rect 155408 197532 155460 197538
rect 155408 197474 155460 197480
rect 155316 191412 155368 191418
rect 155316 191354 155368 191360
rect 155420 191078 155448 197474
rect 155512 196602 155540 197628
rect 155604 196790 155632 199736
rect 155926 199764 155954 200124
rect 155684 199718 155736 199724
rect 155774 199744 155830 199753
rect 155696 196790 155724 199718
rect 155774 199679 155830 199688
rect 155880 199736 155954 199764
rect 156018 199764 156046 200124
rect 156110 199918 156138 200124
rect 156202 199918 156230 200124
rect 156294 199918 156322 200124
rect 156386 199918 156414 200124
rect 156098 199912 156150 199918
rect 156098 199854 156150 199860
rect 156190 199912 156242 199918
rect 156190 199854 156242 199860
rect 156282 199912 156334 199918
rect 156282 199854 156334 199860
rect 156374 199912 156426 199918
rect 156374 199854 156426 199860
rect 156478 199764 156506 200124
rect 156570 199923 156598 200124
rect 156556 199914 156612 199923
rect 156662 199918 156690 200124
rect 156754 199918 156782 200124
rect 156846 199918 156874 200124
rect 156556 199849 156612 199858
rect 156650 199912 156702 199918
rect 156650 199854 156702 199860
rect 156742 199912 156794 199918
rect 156742 199854 156794 199860
rect 156834 199912 156886 199918
rect 156834 199854 156886 199860
rect 156938 199850 156966 200124
rect 157030 199889 157058 200124
rect 157122 199918 157150 200124
rect 157214 199923 157242 200124
rect 157110 199912 157162 199918
rect 157016 199880 157072 199889
rect 156926 199844 156978 199850
rect 157110 199854 157162 199860
rect 157200 199914 157256 199923
rect 157200 199849 157256 199858
rect 157016 199815 157072 199824
rect 156926 199786 156978 199792
rect 156018 199736 156092 199764
rect 155592 196784 155644 196790
rect 155592 196726 155644 196732
rect 155684 196784 155736 196790
rect 155684 196726 155736 196732
rect 155512 196574 155724 196602
rect 155788 196586 155816 199679
rect 155880 198422 155908 199736
rect 155960 199640 156012 199646
rect 155960 199582 156012 199588
rect 155868 198416 155920 198422
rect 155868 198358 155920 198364
rect 155972 198150 156000 199582
rect 155960 198144 156012 198150
rect 155960 198086 156012 198092
rect 155868 196784 155920 196790
rect 155868 196726 155920 196732
rect 155592 196512 155644 196518
rect 155592 196454 155644 196460
rect 155408 191072 155460 191078
rect 155408 191014 155460 191020
rect 155604 188290 155632 196454
rect 155592 188284 155644 188290
rect 155592 188226 155644 188232
rect 155132 187808 155184 187814
rect 155132 187750 155184 187756
rect 154856 184476 154908 184482
rect 154856 184418 154908 184424
rect 155696 151814 155724 196574
rect 155776 196580 155828 196586
rect 155776 196522 155828 196528
rect 155880 191185 155908 196726
rect 156064 196518 156092 199736
rect 156432 199736 156506 199764
rect 156788 199776 156840 199782
rect 156602 199744 156658 199753
rect 156236 199708 156288 199714
rect 156236 199650 156288 199656
rect 156328 199708 156380 199714
rect 156328 199650 156380 199656
rect 156144 199640 156196 199646
rect 156144 199582 156196 199588
rect 156156 196790 156184 199582
rect 156248 199442 156276 199650
rect 156236 199436 156288 199442
rect 156236 199378 156288 199384
rect 156236 199300 156288 199306
rect 156236 199242 156288 199248
rect 156144 196784 156196 196790
rect 156144 196726 156196 196732
rect 156248 196602 156276 199242
rect 156156 196574 156276 196602
rect 156052 196512 156104 196518
rect 156052 196454 156104 196460
rect 156052 195968 156104 195974
rect 156052 195910 156104 195916
rect 155866 191176 155922 191185
rect 155866 191111 155922 191120
rect 155868 191072 155920 191078
rect 155868 191014 155920 191020
rect 155696 151786 155816 151814
rect 154764 151156 154816 151162
rect 154764 151098 154816 151104
rect 155684 142996 155736 143002
rect 155684 142938 155736 142944
rect 154672 140140 154724 140146
rect 154672 140082 154724 140088
rect 155696 139890 155724 142938
rect 155788 140078 155816 151786
rect 155880 144294 155908 191014
rect 156064 151094 156092 195910
rect 156156 181762 156184 196574
rect 156234 196480 156290 196489
rect 156234 196415 156290 196424
rect 156248 183394 156276 196415
rect 156236 183388 156288 183394
rect 156236 183330 156288 183336
rect 156340 182986 156368 199650
rect 156432 196994 156460 199736
rect 156602 199679 156658 199688
rect 156786 199744 156788 199753
rect 157306 199764 157334 200124
rect 157398 199918 157426 200124
rect 157386 199912 157438 199918
rect 157386 199854 157438 199860
rect 157490 199764 157518 200124
rect 156840 199744 156842 199753
rect 157168 199736 157334 199764
rect 157444 199736 157518 199764
rect 156786 199679 156842 199688
rect 157064 199708 157116 199714
rect 156512 199640 156564 199646
rect 156512 199582 156564 199588
rect 156420 196988 156472 196994
rect 156420 196930 156472 196936
rect 156524 196761 156552 199582
rect 156510 196752 156566 196761
rect 156510 196687 156566 196696
rect 156616 196314 156644 199679
rect 157064 199650 157116 199656
rect 156696 199640 156748 199646
rect 156696 199582 156748 199588
rect 156972 199640 157024 199646
rect 156972 199582 157024 199588
rect 156604 196308 156656 196314
rect 156604 196250 156656 196256
rect 156418 196072 156474 196081
rect 156418 196007 156474 196016
rect 156432 189786 156460 196007
rect 156708 190126 156736 199582
rect 156880 199572 156932 199578
rect 156880 199514 156932 199520
rect 156892 198354 156920 199514
rect 156984 199306 157012 199582
rect 156972 199300 157024 199306
rect 156972 199242 157024 199248
rect 156880 198348 156932 198354
rect 156880 198290 156932 198296
rect 156788 196784 156840 196790
rect 156788 196726 156840 196732
rect 156800 192506 156828 196726
rect 156880 196512 156932 196518
rect 156880 196454 156932 196460
rect 156788 192500 156840 192506
rect 156788 192442 156840 192448
rect 156696 190120 156748 190126
rect 156696 190062 156748 190068
rect 156420 189780 156472 189786
rect 156420 189722 156472 189728
rect 156892 188562 156920 196454
rect 156972 196308 157024 196314
rect 156972 196250 157024 196256
rect 156880 188556 156932 188562
rect 156880 188498 156932 188504
rect 156328 182980 156380 182986
rect 156328 182922 156380 182928
rect 156144 181756 156196 181762
rect 156144 181698 156196 181704
rect 156052 151088 156104 151094
rect 156052 151030 156104 151036
rect 155868 144288 155920 144294
rect 155868 144230 155920 144236
rect 156512 141840 156564 141846
rect 156512 141782 156564 141788
rect 155776 140072 155828 140078
rect 155776 140014 155828 140020
rect 156524 139890 156552 141782
rect 156984 141710 157012 196250
rect 157076 195974 157104 199650
rect 157168 199617 157196 199736
rect 157340 199640 157392 199646
rect 157154 199608 157210 199617
rect 157340 199582 157392 199588
rect 157154 199543 157210 199552
rect 157156 199436 157208 199442
rect 157156 199378 157208 199384
rect 157168 197742 157196 199378
rect 157352 199374 157380 199582
rect 157340 199368 157392 199374
rect 157340 199310 157392 199316
rect 157248 199300 157300 199306
rect 157248 199242 157300 199248
rect 157260 198898 157288 199242
rect 157248 198892 157300 198898
rect 157248 198834 157300 198840
rect 157156 197736 157208 197742
rect 157156 197678 157208 197684
rect 157248 196920 157300 196926
rect 157248 196862 157300 196868
rect 157064 195968 157116 195974
rect 157064 195910 157116 195916
rect 157260 195566 157288 196862
rect 157248 195560 157300 195566
rect 157248 195502 157300 195508
rect 157260 189854 157288 195502
rect 157444 194546 157472 199736
rect 157582 199696 157610 200124
rect 157674 199764 157702 200124
rect 157766 199918 157794 200124
rect 157754 199912 157806 199918
rect 157754 199854 157806 199860
rect 157858 199764 157886 200124
rect 157950 199918 157978 200124
rect 158042 199918 158070 200124
rect 158134 199918 158162 200124
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158030 199912 158082 199918
rect 158030 199854 158082 199860
rect 158122 199912 158174 199918
rect 158122 199854 158174 199860
rect 157674 199736 157748 199764
rect 157858 199753 157932 199764
rect 157858 199744 157946 199753
rect 157858 199736 157890 199744
rect 157536 199668 157610 199696
rect 157720 199696 157748 199736
rect 157720 199668 157840 199696
rect 158226 199730 158254 200124
rect 158318 199923 158346 200124
rect 158304 199914 158360 199923
rect 158410 199918 158438 200124
rect 158502 199918 158530 200124
rect 158304 199849 158360 199858
rect 158398 199912 158450 199918
rect 158398 199854 158450 199860
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 158594 199764 158622 200124
rect 158686 199918 158714 200124
rect 158674 199912 158726 199918
rect 158674 199854 158726 199860
rect 158548 199753 158622 199764
rect 157890 199679 157946 199688
rect 157996 199702 158254 199730
rect 158534 199744 158622 199753
rect 158352 199708 158404 199714
rect 157536 196926 157564 199668
rect 157616 199572 157668 199578
rect 157616 199514 157668 199520
rect 157708 199572 157760 199578
rect 157708 199514 157760 199520
rect 157524 196920 157576 196926
rect 157524 196862 157576 196868
rect 157524 196784 157576 196790
rect 157524 196726 157576 196732
rect 157432 194540 157484 194546
rect 157432 194482 157484 194488
rect 157536 189990 157564 196726
rect 157628 194070 157656 199514
rect 157720 196518 157748 199514
rect 157708 196512 157760 196518
rect 157708 196454 157760 196460
rect 157616 194064 157668 194070
rect 157616 194006 157668 194012
rect 157812 193458 157840 199668
rect 157892 199572 157944 199578
rect 157892 199514 157944 199520
rect 157904 198801 157932 199514
rect 157890 198792 157946 198801
rect 157890 198727 157946 198736
rect 157800 193452 157852 193458
rect 157800 193394 157852 193400
rect 157904 193214 157932 198727
rect 157996 194002 158024 199702
rect 158352 199650 158404 199656
rect 158444 199708 158496 199714
rect 158590 199736 158622 199744
rect 158534 199679 158590 199688
rect 158444 199650 158496 199656
rect 158076 199640 158128 199646
rect 158076 199582 158128 199588
rect 158258 199608 158314 199617
rect 158088 196450 158116 199582
rect 158258 199543 158314 199552
rect 158166 198928 158222 198937
rect 158166 198863 158222 198872
rect 158180 196858 158208 198863
rect 158272 196858 158300 199543
rect 158168 196852 158220 196858
rect 158168 196794 158220 196800
rect 158260 196852 158312 196858
rect 158260 196794 158312 196800
rect 158364 196790 158392 199650
rect 158352 196784 158404 196790
rect 158352 196726 158404 196732
rect 158456 196602 158484 199650
rect 158628 199640 158680 199646
rect 158778 199628 158806 200124
rect 158870 199764 158898 200124
rect 158962 199923 158990 200124
rect 158948 199914 159004 199923
rect 158948 199849 159004 199858
rect 158870 199736 158944 199764
rect 158628 199582 158680 199588
rect 158732 199600 158806 199628
rect 158536 199572 158588 199578
rect 158536 199514 158588 199520
rect 158548 197062 158576 199514
rect 158536 197056 158588 197062
rect 158536 196998 158588 197004
rect 158272 196574 158484 196602
rect 158076 196444 158128 196450
rect 158076 196386 158128 196392
rect 158168 196240 158220 196246
rect 158168 196182 158220 196188
rect 157984 193996 158036 194002
rect 157984 193938 158036 193944
rect 157904 193186 158024 193214
rect 157524 189984 157576 189990
rect 157524 189926 157576 189932
rect 157248 189848 157300 189854
rect 157248 189790 157300 189796
rect 157340 144696 157392 144702
rect 157340 144638 157392 144644
rect 157352 143002 157380 144638
rect 157996 144129 158024 193186
rect 158180 184550 158208 196182
rect 158168 184544 158220 184550
rect 158168 184486 158220 184492
rect 158180 180794 158208 184486
rect 158272 184210 158300 196574
rect 158536 196444 158588 196450
rect 158536 196386 158588 196392
rect 158352 193452 158404 193458
rect 158352 193394 158404 193400
rect 158364 187066 158392 193394
rect 158352 187060 158404 187066
rect 158352 187002 158404 187008
rect 158260 184204 158312 184210
rect 158260 184146 158312 184152
rect 158548 182918 158576 196386
rect 158640 195158 158668 199582
rect 158732 198121 158760 199600
rect 158812 199504 158864 199510
rect 158812 199446 158864 199452
rect 158718 198112 158774 198121
rect 158718 198047 158774 198056
rect 158628 195152 158680 195158
rect 158628 195094 158680 195100
rect 158824 190454 158852 199446
rect 158640 190426 158852 190454
rect 158640 189106 158668 190426
rect 158628 189100 158680 189106
rect 158628 189042 158680 189048
rect 158640 187270 158668 189042
rect 158628 187264 158680 187270
rect 158628 187206 158680 187212
rect 158628 186992 158680 186998
rect 158628 186934 158680 186940
rect 158640 186386 158668 186934
rect 158628 186380 158680 186386
rect 158628 186322 158680 186328
rect 158536 182912 158588 182918
rect 158536 182854 158588 182860
rect 158088 180766 158208 180794
rect 158088 144362 158116 180766
rect 158168 144628 158220 144634
rect 158168 144570 158220 144576
rect 158076 144356 158128 144362
rect 158076 144298 158128 144304
rect 157982 144120 158038 144129
rect 157982 144055 158038 144064
rect 157340 142996 157392 143002
rect 157340 142938 157392 142944
rect 157246 142352 157302 142361
rect 157246 142287 157302 142296
rect 156972 141704 157024 141710
rect 156972 141646 157024 141652
rect 157260 139890 157288 142287
rect 158180 139890 158208 144570
rect 158352 141908 158404 141914
rect 158352 141850 158404 141856
rect 158364 140826 158392 141850
rect 158640 141778 158668 186322
rect 158916 183025 158944 199736
rect 159054 199628 159082 200124
rect 159146 199764 159174 200124
rect 159238 199923 159266 200124
rect 159224 199914 159280 199923
rect 159224 199849 159280 199858
rect 159146 199736 159220 199764
rect 159008 199600 159082 199628
rect 159008 196790 159036 199600
rect 159192 198734 159220 199736
rect 159330 199696 159358 200124
rect 159422 199764 159450 200124
rect 159514 199918 159542 200124
rect 159502 199912 159554 199918
rect 159502 199854 159554 199860
rect 159606 199764 159634 200124
rect 159422 199753 159496 199764
rect 159422 199744 159510 199753
rect 159422 199736 159454 199744
rect 159330 199668 159404 199696
rect 159454 199679 159510 199688
rect 159560 199736 159634 199764
rect 159698 199764 159726 200124
rect 159790 199918 159818 200124
rect 159882 199918 159910 200124
rect 159778 199912 159830 199918
rect 159778 199854 159830 199860
rect 159870 199912 159922 199918
rect 159974 199889 160002 200124
rect 159870 199854 159922 199860
rect 159960 199880 160016 199889
rect 159960 199815 160016 199824
rect 160066 199764 160094 200124
rect 159698 199736 159772 199764
rect 159270 199608 159326 199617
rect 159270 199543 159326 199552
rect 159376 199560 159404 199668
rect 159284 199458 159312 199543
rect 159376 199532 159496 199560
rect 159284 199430 159404 199458
rect 159100 198706 159220 198734
rect 158996 196784 159048 196790
rect 158996 196726 159048 196732
rect 159100 196738 159128 198706
rect 159270 197432 159326 197441
rect 159270 197367 159326 197376
rect 159284 197033 159312 197367
rect 159270 197024 159326 197033
rect 159270 196959 159326 196968
rect 159376 196858 159404 199430
rect 159364 196852 159416 196858
rect 159364 196794 159416 196800
rect 159100 196710 159220 196738
rect 159088 196580 159140 196586
rect 159088 196522 159140 196528
rect 159100 184278 159128 196522
rect 159088 184272 159140 184278
rect 159088 184214 159140 184220
rect 158902 183016 158958 183025
rect 158902 182951 158958 182960
rect 159192 181694 159220 196710
rect 159468 196314 159496 199532
rect 159560 196586 159588 199736
rect 159744 199560 159772 199736
rect 159928 199736 160094 199764
rect 159824 199708 159876 199714
rect 159824 199650 159876 199656
rect 159652 199532 159772 199560
rect 159652 199238 159680 199532
rect 159836 199458 159864 199650
rect 159744 199430 159864 199458
rect 159640 199232 159692 199238
rect 159640 199174 159692 199180
rect 159744 198642 159772 199430
rect 159652 198614 159772 198642
rect 159652 197248 159680 198614
rect 159732 198552 159784 198558
rect 159730 198520 159732 198529
rect 159784 198520 159786 198529
rect 159730 198455 159786 198464
rect 159822 198248 159878 198257
rect 159822 198183 159878 198192
rect 159652 197220 159772 197248
rect 159640 197056 159692 197062
rect 159640 196998 159692 197004
rect 159548 196580 159600 196586
rect 159548 196522 159600 196528
rect 159456 196308 159508 196314
rect 159456 196250 159508 196256
rect 159652 191486 159680 196998
rect 159744 196246 159772 197220
rect 159732 196240 159784 196246
rect 159732 196182 159784 196188
rect 159640 191480 159692 191486
rect 159640 191422 159692 191428
rect 159836 183054 159864 198183
rect 159928 191146 159956 199736
rect 160158 199730 160186 200124
rect 160250 199923 160278 200124
rect 160236 199914 160292 199923
rect 160236 199849 160292 199858
rect 160342 199850 160370 200124
rect 160330 199844 160382 199850
rect 160330 199786 160382 199792
rect 160434 199782 160462 200124
rect 160526 199918 160554 200124
rect 160618 199923 160646 200124
rect 160514 199912 160566 199918
rect 160514 199854 160566 199860
rect 160604 199914 160660 199923
rect 160710 199918 160738 200124
rect 160802 199918 160830 200124
rect 160604 199849 160660 199858
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160790 199912 160842 199918
rect 160790 199854 160842 199860
rect 160422 199776 160474 199782
rect 160158 199702 160232 199730
rect 160894 199764 160922 200124
rect 160986 199918 161014 200124
rect 160974 199912 161026 199918
rect 160974 199854 161026 199860
rect 161078 199764 161106 200124
rect 161170 199918 161198 200124
rect 161262 199923 161290 200124
rect 161158 199912 161210 199918
rect 161158 199854 161210 199860
rect 161248 199914 161304 199923
rect 161354 199918 161382 200124
rect 161446 199918 161474 200124
rect 161538 199918 161566 200124
rect 161630 199918 161658 200124
rect 161722 199918 161750 200124
rect 161248 199849 161304 199858
rect 161342 199912 161394 199918
rect 161342 199854 161394 199860
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161526 199912 161578 199918
rect 161526 199854 161578 199860
rect 161618 199912 161670 199918
rect 161618 199854 161670 199860
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161296 199776 161348 199782
rect 160422 199718 160474 199724
rect 160558 199744 160614 199753
rect 160100 199640 160152 199646
rect 160100 199582 160152 199588
rect 160112 199102 160140 199582
rect 160100 199096 160152 199102
rect 160100 199038 160152 199044
rect 160008 196784 160060 196790
rect 160008 196726 160060 196732
rect 160204 196738 160232 199702
rect 160284 199708 160336 199714
rect 160894 199736 160968 199764
rect 161078 199736 161152 199764
rect 160558 199679 160614 199688
rect 160284 199650 160336 199656
rect 160296 197810 160324 199650
rect 160376 199640 160428 199646
rect 160376 199582 160428 199588
rect 160572 199594 160600 199679
rect 160836 199640 160888 199646
rect 160742 199608 160798 199617
rect 160284 197804 160336 197810
rect 160284 197746 160336 197752
rect 159916 191140 159968 191146
rect 159916 191082 159968 191088
rect 160020 186386 160048 196726
rect 160204 196710 160324 196738
rect 160192 196580 160244 196586
rect 160192 196522 160244 196528
rect 160008 186380 160060 186386
rect 160008 186322 160060 186328
rect 159824 183048 159876 183054
rect 159824 182990 159876 182996
rect 159180 181688 159232 181694
rect 159180 181630 159232 181636
rect 160204 144498 160232 196522
rect 160296 144566 160324 196710
rect 160388 196586 160416 199582
rect 160468 199572 160520 199578
rect 160572 199566 160692 199594
rect 160468 199514 160520 199520
rect 160376 196580 160428 196586
rect 160376 196522 160428 196528
rect 160480 196466 160508 199514
rect 160560 199504 160612 199510
rect 160560 199446 160612 199452
rect 160388 196438 160508 196466
rect 160388 149054 160416 196438
rect 160468 195968 160520 195974
rect 160468 195910 160520 195916
rect 160480 184142 160508 195910
rect 160572 185570 160600 199446
rect 160664 190058 160692 199566
rect 160836 199582 160888 199588
rect 160742 199543 160798 199552
rect 160756 199442 160784 199543
rect 160744 199436 160796 199442
rect 160744 199378 160796 199384
rect 160848 198898 160876 199582
rect 160836 198892 160888 198898
rect 160836 198834 160888 198840
rect 160940 198393 160968 199736
rect 161020 199572 161072 199578
rect 161020 199514 161072 199520
rect 160926 198384 160982 198393
rect 160926 198319 160982 198328
rect 160834 197840 160890 197849
rect 160834 197775 160890 197784
rect 160848 197538 160876 197775
rect 160836 197532 160888 197538
rect 160836 197474 160888 197480
rect 160836 196512 160888 196518
rect 160836 196454 160888 196460
rect 160848 192574 160876 196454
rect 160836 192568 160888 192574
rect 160836 192510 160888 192516
rect 161032 190454 161060 199514
rect 161124 198490 161152 199736
rect 161572 199776 161624 199782
rect 161296 199718 161348 199724
rect 161478 199744 161534 199753
rect 161204 199708 161256 199714
rect 161204 199650 161256 199656
rect 161112 198484 161164 198490
rect 161112 198426 161164 198432
rect 161216 196761 161244 199650
rect 161202 196752 161258 196761
rect 161202 196687 161258 196696
rect 161308 195974 161336 199718
rect 161572 199718 161624 199724
rect 161662 199744 161718 199753
rect 161478 199679 161534 199688
rect 161388 199640 161440 199646
rect 161388 199582 161440 199588
rect 161400 197266 161428 199582
rect 161388 197260 161440 197266
rect 161388 197202 161440 197208
rect 161492 197130 161520 199679
rect 161480 197124 161532 197130
rect 161480 197066 161532 197072
rect 161480 196240 161532 196246
rect 161480 196182 161532 196188
rect 161296 195968 161348 195974
rect 161296 195910 161348 195916
rect 161032 190426 161336 190454
rect 160652 190052 160704 190058
rect 160652 189994 160704 190000
rect 160560 185564 160612 185570
rect 160560 185506 160612 185512
rect 160468 184136 160520 184142
rect 160468 184078 160520 184084
rect 160376 149048 160428 149054
rect 160376 148990 160428 148996
rect 160376 145784 160428 145790
rect 160376 145726 160428 145732
rect 160284 144560 160336 144566
rect 160284 144502 160336 144508
rect 160192 144492 160244 144498
rect 160192 144434 160244 144440
rect 159824 142996 159876 143002
rect 159824 142938 159876 142944
rect 158628 141772 158680 141778
rect 158628 141714 158680 141720
rect 158352 140820 158404 140826
rect 158352 140762 158404 140768
rect 154500 139862 154560 139890
rect 155388 139862 155724 139890
rect 156216 139862 156552 139890
rect 157044 139862 157288 139890
rect 157872 139862 158208 139890
rect 158364 139890 158392 140762
rect 159836 139890 159864 142938
rect 160388 140162 160416 145726
rect 161308 144430 161336 190426
rect 161492 185502 161520 196182
rect 161480 185496 161532 185502
rect 161480 185438 161532 185444
rect 161584 148714 161612 199718
rect 161814 199730 161842 200124
rect 161906 199918 161934 200124
rect 161998 199918 162026 200124
rect 162090 199918 162118 200124
rect 161894 199912 161946 199918
rect 161894 199854 161946 199860
rect 161986 199912 162038 199918
rect 161986 199854 162038 199860
rect 162078 199912 162130 199918
rect 162078 199854 162130 199860
rect 161814 199702 161888 199730
rect 161662 199679 161718 199688
rect 161676 196450 161704 199679
rect 161756 199640 161808 199646
rect 161756 199582 161808 199588
rect 161664 196444 161716 196450
rect 161664 196386 161716 196392
rect 161664 196104 161716 196110
rect 161664 196046 161716 196052
rect 161676 178770 161704 196046
rect 161768 195294 161796 199582
rect 161860 197674 161888 199702
rect 162182 199696 162210 200124
rect 162274 199918 162302 200124
rect 162262 199912 162314 199918
rect 162262 199854 162314 199860
rect 162366 199764 162394 200124
rect 162136 199668 162210 199696
rect 162320 199736 162394 199764
rect 162032 199640 162084 199646
rect 162032 199582 162084 199588
rect 161940 199504 161992 199510
rect 161940 199446 161992 199452
rect 161952 198665 161980 199446
rect 161938 198656 161994 198665
rect 161938 198591 161994 198600
rect 161940 198484 161992 198490
rect 161940 198426 161992 198432
rect 161848 197668 161900 197674
rect 161848 197610 161900 197616
rect 161756 195288 161808 195294
rect 161756 195230 161808 195236
rect 161952 191554 161980 198426
rect 162044 197441 162072 199582
rect 162030 197432 162086 197441
rect 162030 197367 162086 197376
rect 161940 191548 161992 191554
rect 161940 191490 161992 191496
rect 162136 191434 162164 199668
rect 162216 199436 162268 199442
rect 162216 199378 162268 199384
rect 161768 191406 162164 191434
rect 161768 185910 161796 191406
rect 162228 186998 162256 199378
rect 162320 193214 162348 199736
rect 162458 199696 162486 200124
rect 162550 199764 162578 200124
rect 162642 199889 162670 200124
rect 162628 199880 162684 199889
rect 162628 199815 162684 199824
rect 162734 199764 162762 200124
rect 162550 199736 162624 199764
rect 162412 199668 162486 199696
rect 162412 196110 162440 199668
rect 162492 199572 162544 199578
rect 162492 199514 162544 199520
rect 162504 199345 162532 199514
rect 162490 199336 162546 199345
rect 162490 199271 162546 199280
rect 162400 196104 162452 196110
rect 162400 196046 162452 196052
rect 162596 193934 162624 199736
rect 162688 199736 162762 199764
rect 162826 199764 162854 200124
rect 162918 199918 162946 200124
rect 162906 199912 162958 199918
rect 162906 199854 162958 199860
rect 163010 199764 163038 200124
rect 163102 199918 163130 200124
rect 163194 199918 163222 200124
rect 163286 199918 163314 200124
rect 163090 199912 163142 199918
rect 163090 199854 163142 199860
rect 163182 199912 163234 199918
rect 163182 199854 163234 199860
rect 163274 199912 163326 199918
rect 163274 199854 163326 199860
rect 162826 199736 162900 199764
rect 162688 196246 162716 199736
rect 162768 199640 162820 199646
rect 162768 199582 162820 199588
rect 162780 198082 162808 199582
rect 162872 198490 162900 199736
rect 162964 199736 163038 199764
rect 162860 198484 162912 198490
rect 162860 198426 162912 198432
rect 162768 198076 162820 198082
rect 162768 198018 162820 198024
rect 162676 196240 162728 196246
rect 162676 196182 162728 196188
rect 162584 193928 162636 193934
rect 162584 193870 162636 193876
rect 162320 193186 162440 193214
rect 162216 186992 162268 186998
rect 162216 186934 162268 186940
rect 161756 185904 161808 185910
rect 161756 185846 161808 185852
rect 161664 178764 161716 178770
rect 161664 178706 161716 178712
rect 162412 151814 162440 193186
rect 162676 191548 162728 191554
rect 162676 191490 162728 191496
rect 162688 191350 162716 191490
rect 162676 191344 162728 191350
rect 162676 191286 162728 191292
rect 162676 185904 162728 185910
rect 162676 185846 162728 185852
rect 162688 182102 162716 185846
rect 162676 182096 162728 182102
rect 162676 182038 162728 182044
rect 162412 151786 162532 151814
rect 161572 148708 161624 148714
rect 161572 148650 161624 148656
rect 162400 145648 162452 145654
rect 162400 145590 162452 145596
rect 161296 144424 161348 144430
rect 161296 144366 161348 144372
rect 162308 143064 162360 143070
rect 162308 143006 162360 143012
rect 161388 142180 161440 142186
rect 161388 142122 161440 142128
rect 158364 139862 158700 139890
rect 159528 139862 159864 139890
rect 160342 140134 160416 140162
rect 160342 139876 160370 140134
rect 161400 139890 161428 142122
rect 162320 139890 162348 143006
rect 161184 139862 161428 139890
rect 162012 139862 162348 139890
rect 162412 139890 162440 145590
rect 162504 145586 162532 151786
rect 162492 145580 162544 145586
rect 162492 145522 162544 145528
rect 162780 140185 162808 198018
rect 162964 197946 162992 199736
rect 163044 199640 163096 199646
rect 163378 199628 163406 200124
rect 163470 199764 163498 200124
rect 163562 199889 163590 200124
rect 163548 199880 163604 199889
rect 163548 199815 163604 199824
rect 163654 199764 163682 200124
rect 163746 199918 163774 200124
rect 163734 199912 163786 199918
rect 163734 199854 163786 199860
rect 163470 199736 163544 199764
rect 163654 199736 163728 199764
rect 163332 199600 163406 199628
rect 163096 199588 163176 199594
rect 163044 199582 163176 199588
rect 163056 199566 163176 199582
rect 163044 199504 163096 199510
rect 163044 199446 163096 199452
rect 162952 197940 163004 197946
rect 162952 197882 163004 197888
rect 162952 196444 163004 196450
rect 162952 196386 163004 196392
rect 162964 145994 162992 196386
rect 163056 148850 163084 199446
rect 163148 196790 163176 199566
rect 163228 199572 163280 199578
rect 163228 199514 163280 199520
rect 163240 197985 163268 199514
rect 163226 197976 163282 197985
rect 163226 197911 163282 197920
rect 163226 197840 163282 197849
rect 163226 197775 163282 197784
rect 163136 196784 163188 196790
rect 163136 196726 163188 196732
rect 163240 196602 163268 197775
rect 163148 196574 163268 196602
rect 163148 153882 163176 196574
rect 163332 195974 163360 199600
rect 163516 197033 163544 199736
rect 163596 198892 163648 198898
rect 163596 198834 163648 198840
rect 163608 198626 163636 198834
rect 163596 198620 163648 198626
rect 163596 198562 163648 198568
rect 163502 197024 163558 197033
rect 163502 196959 163558 196968
rect 163504 196852 163556 196858
rect 163504 196794 163556 196800
rect 163320 195968 163372 195974
rect 163320 195910 163372 195916
rect 163228 194540 163280 194546
rect 163228 194482 163280 194488
rect 163240 188426 163268 194482
rect 163516 190194 163544 196794
rect 163700 196761 163728 199736
rect 163838 199696 163866 200124
rect 163930 199764 163958 200124
rect 164022 199889 164050 200124
rect 164008 199880 164064 199889
rect 164114 199850 164142 200124
rect 164206 199918 164234 200124
rect 164194 199912 164246 199918
rect 164194 199854 164246 199860
rect 164008 199815 164064 199824
rect 164102 199844 164154 199850
rect 164102 199786 164154 199792
rect 163930 199736 164004 199764
rect 163838 199668 163912 199696
rect 163780 199504 163832 199510
rect 163780 199446 163832 199452
rect 163686 196752 163742 196761
rect 163686 196687 163742 196696
rect 163688 196580 163740 196586
rect 163688 196522 163740 196528
rect 163700 192914 163728 196522
rect 163688 192908 163740 192914
rect 163688 192850 163740 192856
rect 163504 190188 163556 190194
rect 163504 190130 163556 190136
rect 163594 189136 163650 189145
rect 163594 189071 163650 189080
rect 163228 188420 163280 188426
rect 163228 188362 163280 188368
rect 163608 187542 163636 189071
rect 163596 187536 163648 187542
rect 163596 187478 163648 187484
rect 163700 187338 163728 192850
rect 163688 187332 163740 187338
rect 163688 187274 163740 187280
rect 163136 153876 163188 153882
rect 163136 153818 163188 153824
rect 163044 148844 163096 148850
rect 163044 148786 163096 148792
rect 162952 145988 163004 145994
rect 162952 145930 163004 145936
rect 163792 140282 163820 199446
rect 163884 194546 163912 199668
rect 163976 199510 164004 199736
rect 164056 199708 164108 199714
rect 164056 199650 164108 199656
rect 164148 199708 164200 199714
rect 164148 199650 164200 199656
rect 163964 199504 164016 199510
rect 163964 199446 164016 199452
rect 164068 199050 164096 199650
rect 163976 199022 164096 199050
rect 163976 196450 164004 199022
rect 164056 198960 164108 198966
rect 164054 198928 164056 198937
rect 164108 198928 164110 198937
rect 164054 198863 164110 198872
rect 164056 197260 164108 197266
rect 164056 197202 164108 197208
rect 164068 196518 164096 197202
rect 164160 196586 164188 199650
rect 164298 199628 164326 200124
rect 164390 199730 164418 200124
rect 164482 199918 164510 200124
rect 164470 199912 164522 199918
rect 164470 199854 164522 199860
rect 164390 199702 164464 199730
rect 164298 199600 164372 199628
rect 164240 199504 164292 199510
rect 164240 199446 164292 199452
rect 164252 198966 164280 199446
rect 164240 198960 164292 198966
rect 164240 198902 164292 198908
rect 164344 198529 164372 199600
rect 164330 198520 164386 198529
rect 164330 198455 164386 198464
rect 164240 198212 164292 198218
rect 164240 198154 164292 198160
rect 164252 197985 164280 198154
rect 164238 197976 164294 197985
rect 164238 197911 164294 197920
rect 164240 197736 164292 197742
rect 164240 197678 164292 197684
rect 164252 196625 164280 197678
rect 164238 196616 164294 196625
rect 164148 196580 164200 196586
rect 164238 196551 164294 196560
rect 164148 196522 164200 196528
rect 164056 196512 164108 196518
rect 164056 196454 164108 196460
rect 164436 196450 164464 199702
rect 164574 199696 164602 200124
rect 164666 199918 164694 200124
rect 164758 199918 164786 200124
rect 164850 199918 164878 200124
rect 164942 199918 164970 200124
rect 164654 199912 164706 199918
rect 164654 199854 164706 199860
rect 164746 199912 164798 199918
rect 164746 199854 164798 199860
rect 164838 199912 164890 199918
rect 164838 199854 164890 199860
rect 164930 199912 164982 199918
rect 164930 199854 164982 199860
rect 165034 199764 165062 200124
rect 165126 199918 165154 200124
rect 165218 199923 165246 200124
rect 165114 199912 165166 199918
rect 165114 199854 165166 199860
rect 165204 199914 165260 199923
rect 165204 199849 165260 199858
rect 164988 199736 165062 199764
rect 165158 199744 165214 199753
rect 164528 199668 164602 199696
rect 164884 199708 164936 199714
rect 164528 199617 164556 199668
rect 164884 199650 164936 199656
rect 164896 199617 164924 199650
rect 164514 199608 164570 199617
rect 164882 199608 164938 199617
rect 164514 199543 164570 199552
rect 164700 199572 164752 199578
rect 164882 199543 164938 199552
rect 164700 199514 164752 199520
rect 164516 199504 164568 199510
rect 164516 199446 164568 199452
rect 164608 199504 164660 199510
rect 164608 199446 164660 199452
rect 163964 196444 164016 196450
rect 163964 196386 164016 196392
rect 164424 196444 164476 196450
rect 164424 196386 164476 196392
rect 164528 195956 164556 199446
rect 164620 196568 164648 199446
rect 164712 196761 164740 199514
rect 164884 199504 164936 199510
rect 164884 199446 164936 199452
rect 164792 198960 164844 198966
rect 164896 198937 164924 199446
rect 164792 198902 164844 198908
rect 164882 198928 164938 198937
rect 164804 198665 164832 198902
rect 164882 198863 164938 198872
rect 164790 198656 164846 198665
rect 164790 198591 164846 198600
rect 164896 197354 164924 198863
rect 164988 197470 165016 199736
rect 165310 199730 165338 200124
rect 165214 199702 165338 199730
rect 165158 199679 165214 199688
rect 165068 199640 165120 199646
rect 165402 199628 165430 200124
rect 165494 199696 165522 200124
rect 165586 199764 165614 200124
rect 165678 199889 165706 200124
rect 165664 199880 165720 199889
rect 165664 199815 165720 199824
rect 165586 199736 165660 199764
rect 165494 199668 165568 199696
rect 165068 199582 165120 199588
rect 165356 199600 165430 199628
rect 164976 197464 165028 197470
rect 164976 197406 165028 197412
rect 164896 197326 165016 197354
rect 164698 196752 164754 196761
rect 164698 196687 164754 196696
rect 164620 196540 164832 196568
rect 164700 196444 164752 196450
rect 164700 196386 164752 196392
rect 164436 195928 164556 195956
rect 163872 194540 163924 194546
rect 163872 194482 163924 194488
rect 164148 187536 164200 187542
rect 164148 187478 164200 187484
rect 164160 186930 164188 187478
rect 164148 186924 164200 186930
rect 164148 186866 164200 186872
rect 164436 178702 164464 195928
rect 164514 195392 164570 195401
rect 164514 195327 164570 195336
rect 164528 183122 164556 195327
rect 164608 195084 164660 195090
rect 164608 195026 164660 195032
rect 164620 184686 164648 195026
rect 164712 185842 164740 196386
rect 164804 194478 164832 196540
rect 164884 195424 164936 195430
rect 164884 195366 164936 195372
rect 164792 194472 164844 194478
rect 164792 194414 164844 194420
rect 164896 193526 164924 195366
rect 164988 193526 165016 197326
rect 165080 194886 165108 199582
rect 165252 199436 165304 199442
rect 165252 199378 165304 199384
rect 165158 198792 165214 198801
rect 165158 198727 165214 198736
rect 165172 195430 165200 198727
rect 165160 195424 165212 195430
rect 165160 195366 165212 195372
rect 165160 195288 165212 195294
rect 165160 195230 165212 195236
rect 165068 194880 165120 194886
rect 165068 194822 165120 194828
rect 164884 193520 164936 193526
rect 164884 193462 164936 193468
rect 164976 193520 165028 193526
rect 164976 193462 165028 193468
rect 164700 185836 164752 185842
rect 164700 185778 164752 185784
rect 164608 184680 164660 184686
rect 164608 184622 164660 184628
rect 164896 184482 164924 193462
rect 164884 184476 164936 184482
rect 164884 184418 164936 184424
rect 164516 183116 164568 183122
rect 164516 183058 164568 183064
rect 164424 178696 164476 178702
rect 164424 178638 164476 178644
rect 164332 145716 164384 145722
rect 164332 145658 164384 145664
rect 163872 143132 163924 143138
rect 163872 143074 163924 143080
rect 163780 140276 163832 140282
rect 163780 140218 163832 140224
rect 162766 140176 162822 140185
rect 162766 140111 162822 140120
rect 163884 139890 163912 143074
rect 164344 140758 164372 145658
rect 164422 145616 164478 145625
rect 164422 145551 164478 145560
rect 164332 140752 164384 140758
rect 164332 140694 164384 140700
rect 162412 139862 162840 139890
rect 163668 139862 163912 139890
rect 164436 139890 164464 145551
rect 165172 141574 165200 195230
rect 165264 148918 165292 199378
rect 165356 195294 165384 199600
rect 165436 199368 165488 199374
rect 165436 199310 165488 199316
rect 165448 198898 165476 199310
rect 165436 198892 165488 198898
rect 165436 198834 165488 198840
rect 165434 198792 165490 198801
rect 165434 198727 165436 198736
rect 165488 198727 165490 198736
rect 165436 198698 165488 198704
rect 165436 198416 165488 198422
rect 165436 198358 165488 198364
rect 165448 198082 165476 198358
rect 165436 198076 165488 198082
rect 165436 198018 165488 198024
rect 165434 197976 165490 197985
rect 165434 197911 165490 197920
rect 165448 195702 165476 197911
rect 165436 195696 165488 195702
rect 165436 195638 165488 195644
rect 165344 195288 165396 195294
rect 165344 195230 165396 195236
rect 165434 195256 165490 195265
rect 165434 195191 165490 195200
rect 165448 194970 165476 195191
rect 165540 195090 165568 199668
rect 165632 198694 165660 199736
rect 165770 199696 165798 200124
rect 165862 199918 165890 200124
rect 165954 199918 165982 200124
rect 165850 199912 165902 199918
rect 165850 199854 165902 199860
rect 165942 199912 165994 199918
rect 166046 199889 166074 200124
rect 166138 199918 166166 200124
rect 166126 199912 166178 199918
rect 165942 199854 165994 199860
rect 166032 199880 166088 199889
rect 166230 199889 166258 200124
rect 166126 199854 166178 199860
rect 166216 199880 166272 199889
rect 166032 199815 166088 199824
rect 166322 199850 166350 200124
rect 166216 199815 166272 199824
rect 166310 199844 166362 199850
rect 166310 199786 166362 199792
rect 166080 199776 166132 199782
rect 166080 199718 166132 199724
rect 165988 199708 166040 199714
rect 165770 199668 165844 199696
rect 165620 198688 165672 198694
rect 165620 198630 165672 198636
rect 165712 198348 165764 198354
rect 165712 198290 165764 198296
rect 165620 197532 165672 197538
rect 165620 197474 165672 197480
rect 165528 195084 165580 195090
rect 165528 195026 165580 195032
rect 165448 194942 165568 194970
rect 165436 194880 165488 194886
rect 165436 194822 165488 194828
rect 165448 191690 165476 194822
rect 165436 191684 165488 191690
rect 165436 191626 165488 191632
rect 165448 184414 165476 191626
rect 165540 187202 165568 194942
rect 165632 193730 165660 197474
rect 165724 195566 165752 198290
rect 165712 195560 165764 195566
rect 165712 195502 165764 195508
rect 165712 195424 165764 195430
rect 165712 195366 165764 195372
rect 165620 193724 165672 193730
rect 165620 193666 165672 193672
rect 165620 193520 165672 193526
rect 165620 193462 165672 193468
rect 165528 187196 165580 187202
rect 165528 187138 165580 187144
rect 165528 184680 165580 184686
rect 165528 184622 165580 184628
rect 165436 184408 165488 184414
rect 165436 184350 165488 184356
rect 165540 184346 165568 184622
rect 165528 184340 165580 184346
rect 165528 184282 165580 184288
rect 165252 148912 165304 148918
rect 165252 148854 165304 148860
rect 165632 141817 165660 193462
rect 165724 147082 165752 195366
rect 165816 147150 165844 199668
rect 165988 199650 166040 199656
rect 165896 199436 165948 199442
rect 165896 199378 165948 199384
rect 165908 199345 165936 199378
rect 165894 199336 165950 199345
rect 165894 199271 165950 199280
rect 165896 198416 165948 198422
rect 165896 198358 165948 198364
rect 165908 197441 165936 198358
rect 165894 197432 165950 197441
rect 165894 197367 165950 197376
rect 166000 196636 166028 199650
rect 166092 197062 166120 199718
rect 166264 199708 166316 199714
rect 166264 199650 166316 199656
rect 166172 198892 166224 198898
rect 166172 198834 166224 198840
rect 166080 197056 166132 197062
rect 166080 196998 166132 197004
rect 166000 196608 166120 196636
rect 165988 196444 166040 196450
rect 165988 196386 166040 196392
rect 165896 195288 165948 195294
rect 165896 195230 165948 195236
rect 165908 151230 165936 195230
rect 166000 183190 166028 196386
rect 166092 187406 166120 196608
rect 166184 196178 166212 198834
rect 166276 198490 166304 199650
rect 166414 199628 166442 200124
rect 166506 199764 166534 200124
rect 166598 199889 166626 200124
rect 166690 199918 166718 200124
rect 166782 199918 166810 200124
rect 166874 199923 166902 200124
rect 166678 199912 166730 199918
rect 166584 199880 166640 199889
rect 166678 199854 166730 199860
rect 166770 199912 166822 199918
rect 166770 199854 166822 199860
rect 166860 199914 166916 199923
rect 166860 199849 166916 199858
rect 166584 199815 166640 199824
rect 166724 199776 166776 199782
rect 166506 199736 166580 199764
rect 166368 199600 166442 199628
rect 166264 198484 166316 198490
rect 166264 198426 166316 198432
rect 166172 196172 166224 196178
rect 166172 196114 166224 196120
rect 166368 195634 166396 199600
rect 166552 195650 166580 199736
rect 166724 199718 166776 199724
rect 166814 199744 166870 199753
rect 166632 199368 166684 199374
rect 166632 199310 166684 199316
rect 166356 195628 166408 195634
rect 166356 195570 166408 195576
rect 166460 195622 166580 195650
rect 166460 195430 166488 195622
rect 166540 195560 166592 195566
rect 166540 195502 166592 195508
rect 166448 195424 166500 195430
rect 166448 195366 166500 195372
rect 166552 194818 166580 195502
rect 166540 194812 166592 194818
rect 166540 194754 166592 194760
rect 166644 187610 166672 199310
rect 166736 195294 166764 199718
rect 166814 199679 166870 199688
rect 166828 196450 166856 199679
rect 166966 199594 166994 200124
rect 167058 199850 167086 200124
rect 167150 199918 167178 200124
rect 167242 199918 167270 200124
rect 167334 199923 167362 200124
rect 167138 199912 167190 199918
rect 167138 199854 167190 199860
rect 167230 199912 167282 199918
rect 167230 199854 167282 199860
rect 167320 199914 167376 199923
rect 167426 199918 167454 200124
rect 167518 199923 167546 200124
rect 167046 199844 167098 199850
rect 167320 199849 167376 199858
rect 167414 199912 167466 199918
rect 167414 199854 167466 199860
rect 167504 199914 167560 199923
rect 167504 199849 167560 199858
rect 167046 199786 167098 199792
rect 167458 199744 167514 199753
rect 167092 199708 167144 199714
rect 167610 199696 167638 200124
rect 167702 199764 167730 200124
rect 167794 199918 167822 200124
rect 167886 199918 167914 200124
rect 167978 199918 168006 200124
rect 168070 199918 168098 200124
rect 168162 199918 168190 200124
rect 167782 199912 167834 199918
rect 167782 199854 167834 199860
rect 167874 199912 167926 199918
rect 167874 199854 167926 199860
rect 167966 199912 168018 199918
rect 167966 199854 168018 199860
rect 168058 199912 168110 199918
rect 168058 199854 168110 199860
rect 168150 199912 168202 199918
rect 168150 199854 168202 199860
rect 167702 199736 167776 199764
rect 167458 199679 167514 199688
rect 167092 199650 167144 199656
rect 166966 199566 167040 199594
rect 166816 196444 166868 196450
rect 166816 196386 166868 196392
rect 167012 196382 167040 199566
rect 167104 198393 167132 199650
rect 167276 199572 167328 199578
rect 167276 199514 167328 199520
rect 167184 199436 167236 199442
rect 167184 199378 167236 199384
rect 167090 198384 167146 198393
rect 167090 198319 167146 198328
rect 167000 196376 167052 196382
rect 167000 196318 167052 196324
rect 167000 196104 167052 196110
rect 167000 196046 167052 196052
rect 166724 195288 166776 195294
rect 166724 195230 166776 195236
rect 167012 194274 167040 196046
rect 167000 194268 167052 194274
rect 167000 194210 167052 194216
rect 167012 191214 167040 194210
rect 167000 191208 167052 191214
rect 167000 191150 167052 191156
rect 166632 187604 166684 187610
rect 166632 187546 166684 187552
rect 166080 187400 166132 187406
rect 166080 187342 166132 187348
rect 165988 183184 166040 183190
rect 165988 183126 166040 183132
rect 165896 151224 165948 151230
rect 165896 151166 165948 151172
rect 167196 148306 167224 199378
rect 167288 196654 167316 199514
rect 167368 199368 167420 199374
rect 167368 199310 167420 199316
rect 167276 196648 167328 196654
rect 167276 196590 167328 196596
rect 167380 196110 167408 199310
rect 167368 196104 167420 196110
rect 167368 196046 167420 196052
rect 167368 195288 167420 195294
rect 167368 195230 167420 195236
rect 167276 191004 167328 191010
rect 167276 190946 167328 190952
rect 167288 148782 167316 190946
rect 167380 180198 167408 195230
rect 167472 187474 167500 199679
rect 167564 199668 167638 199696
rect 167564 191010 167592 199668
rect 167644 199572 167696 199578
rect 167644 199514 167696 199520
rect 167656 198937 167684 199514
rect 167642 198928 167698 198937
rect 167642 198863 167698 198872
rect 167644 198756 167696 198762
rect 167644 198698 167696 198704
rect 167656 197713 167684 198698
rect 167642 197704 167698 197713
rect 167642 197639 167698 197648
rect 167552 191004 167604 191010
rect 167552 190946 167604 190952
rect 167748 190454 167776 199736
rect 168254 199730 168282 200124
rect 168346 199918 168374 200124
rect 168438 199918 168466 200124
rect 168334 199912 168386 199918
rect 168334 199854 168386 199860
rect 168426 199912 168478 199918
rect 168426 199854 168478 199860
rect 168530 199764 168558 200124
rect 168622 199889 168650 200124
rect 168608 199880 168664 199889
rect 168608 199815 168664 199824
rect 168714 199764 168742 200124
rect 168484 199736 168558 199764
rect 168668 199736 168742 199764
rect 168254 199702 168328 199730
rect 168012 199572 168064 199578
rect 168012 199514 168064 199520
rect 168104 199572 168156 199578
rect 168104 199514 168156 199520
rect 167920 199504 167972 199510
rect 167920 199446 167972 199452
rect 167932 196858 167960 199446
rect 168024 197554 168052 199514
rect 168116 197713 168144 199514
rect 168102 197704 168158 197713
rect 168102 197639 168158 197648
rect 168024 197526 168144 197554
rect 168012 197464 168064 197470
rect 168012 197406 168064 197412
rect 167920 196852 167972 196858
rect 167920 196794 167972 196800
rect 168024 193905 168052 197406
rect 168116 196466 168144 197526
rect 168116 196438 168236 196466
rect 168102 196344 168158 196353
rect 168102 196279 168158 196288
rect 168010 193896 168066 193905
rect 168010 193831 168066 193840
rect 167748 190426 168052 190454
rect 167460 187468 167512 187474
rect 167460 187410 167512 187416
rect 167644 184748 167696 184754
rect 167644 184690 167696 184696
rect 167368 180192 167420 180198
rect 167368 180134 167420 180140
rect 167656 178838 167684 184690
rect 167644 178832 167696 178838
rect 167644 178774 167696 178780
rect 167276 148776 167328 148782
rect 167276 148718 167328 148724
rect 167184 148300 167236 148306
rect 167184 148242 167236 148248
rect 168024 147218 168052 190426
rect 168116 148646 168144 196279
rect 168208 184754 168236 196438
rect 168300 195294 168328 199702
rect 168380 199708 168432 199714
rect 168380 199650 168432 199656
rect 168392 199050 168420 199650
rect 168484 199510 168512 199736
rect 168564 199640 168616 199646
rect 168668 199617 168696 199736
rect 168806 199696 168834 200124
rect 168760 199668 168834 199696
rect 168564 199582 168616 199588
rect 168654 199608 168710 199617
rect 168472 199504 168524 199510
rect 168472 199446 168524 199452
rect 168392 199022 168512 199050
rect 168378 198928 168434 198937
rect 168378 198863 168434 198872
rect 168392 198762 168420 198863
rect 168380 198756 168432 198762
rect 168380 198698 168432 198704
rect 168484 198354 168512 199022
rect 168472 198348 168524 198354
rect 168472 198290 168524 198296
rect 168576 198234 168604 199582
rect 168654 199543 168710 199552
rect 168656 199436 168708 199442
rect 168656 199378 168708 199384
rect 168392 198206 168604 198234
rect 168288 195288 168340 195294
rect 168288 195230 168340 195236
rect 168196 184748 168248 184754
rect 168196 184690 168248 184696
rect 168104 148640 168156 148646
rect 168104 148582 168156 148588
rect 168012 147212 168064 147218
rect 168012 147154 168064 147160
rect 165804 147144 165856 147150
rect 165804 147086 165856 147092
rect 165712 147076 165764 147082
rect 165712 147018 165764 147024
rect 168392 147014 168420 198206
rect 168668 197402 168696 199378
rect 168656 197396 168708 197402
rect 168656 197338 168708 197344
rect 168760 196636 168788 199668
rect 168898 199560 168926 200124
rect 168668 196608 168788 196636
rect 168852 199532 168926 199560
rect 168472 196580 168524 196586
rect 168472 196522 168524 196528
rect 168484 148481 168512 196522
rect 168564 196444 168616 196450
rect 168564 196386 168616 196392
rect 168576 148578 168604 196386
rect 168668 180130 168696 196608
rect 168748 196240 168800 196246
rect 168748 196182 168800 196188
rect 168760 186402 168788 196182
rect 168852 195566 168880 199532
rect 168990 199492 169018 200124
rect 169082 199918 169110 200124
rect 169070 199912 169122 199918
rect 169070 199854 169122 199860
rect 169174 199764 169202 200124
rect 169266 199889 169294 200124
rect 169358 199918 169386 200124
rect 169346 199912 169398 199918
rect 169252 199880 169308 199889
rect 169450 199889 169478 200124
rect 169346 199854 169398 199860
rect 169436 199880 169492 199889
rect 169252 199815 169308 199824
rect 169436 199815 169492 199824
rect 169300 199776 169352 199782
rect 169174 199736 169248 199764
rect 169116 199640 169168 199646
rect 169116 199582 169168 199588
rect 168944 199464 169018 199492
rect 168944 196450 168972 199464
rect 169128 199186 169156 199582
rect 169036 199158 169156 199186
rect 169036 198286 169064 199158
rect 169220 199050 169248 199736
rect 169300 199718 169352 199724
rect 169312 199458 169340 199718
rect 169542 199696 169570 200124
rect 169634 199918 169662 200124
rect 169622 199912 169674 199918
rect 169622 199854 169674 199860
rect 169726 199730 169754 200124
rect 169818 199918 169846 200124
rect 169910 199923 169938 200124
rect 169806 199912 169858 199918
rect 169806 199854 169858 199860
rect 169896 199914 169952 199923
rect 170002 199918 170030 200124
rect 170094 199918 170122 200124
rect 170186 199918 170214 200124
rect 169896 199849 169952 199858
rect 169990 199912 170042 199918
rect 169990 199854 170042 199860
rect 170082 199912 170134 199918
rect 170082 199854 170134 199860
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 169944 199776 169996 199782
rect 169850 199744 169906 199753
rect 169496 199668 169570 199696
rect 169622 199708 169674 199714
rect 169390 199608 169446 199617
rect 169390 199543 169392 199552
rect 169444 199543 169446 199552
rect 169392 199514 169444 199520
rect 169312 199430 169432 199458
rect 169128 199022 169248 199050
rect 169024 198280 169076 198286
rect 169024 198222 169076 198228
rect 169024 196648 169076 196654
rect 169024 196590 169076 196596
rect 168932 196444 168984 196450
rect 168932 196386 168984 196392
rect 168840 195560 168892 195566
rect 168840 195502 168892 195508
rect 169036 194886 169064 196590
rect 169024 194880 169076 194886
rect 169024 194822 169076 194828
rect 169128 193214 169156 199022
rect 169208 198892 169260 198898
rect 169208 198834 169260 198840
rect 169220 198558 169248 198834
rect 169208 198552 169260 198558
rect 169208 198494 169260 198500
rect 169208 198416 169260 198422
rect 169208 198358 169260 198364
rect 169220 198286 169248 198358
rect 169208 198280 169260 198286
rect 169208 198222 169260 198228
rect 169300 198144 169352 198150
rect 169300 198086 169352 198092
rect 169208 196852 169260 196858
rect 169208 196794 169260 196800
rect 168944 193186 169156 193214
rect 168838 191720 168894 191729
rect 168838 191655 168894 191664
rect 168852 190534 168880 191655
rect 168840 190528 168892 190534
rect 168840 190470 168892 190476
rect 168944 187542 168972 193186
rect 168932 187536 168984 187542
rect 168932 187478 168984 187484
rect 168760 186374 168880 186402
rect 168748 186108 168800 186114
rect 168748 186050 168800 186056
rect 168760 186017 168788 186050
rect 168746 186008 168802 186017
rect 168746 185943 168802 185952
rect 168760 184958 168788 185943
rect 168748 184952 168800 184958
rect 168748 184894 168800 184900
rect 168852 184770 168880 186374
rect 169220 185774 169248 196794
rect 169312 189650 169340 198086
rect 169404 198082 169432 199430
rect 169392 198076 169444 198082
rect 169392 198018 169444 198024
rect 169392 197804 169444 197810
rect 169392 197746 169444 197752
rect 169404 190262 169432 197746
rect 169496 196586 169524 199668
rect 169726 199702 169800 199730
rect 169622 199650 169674 199656
rect 169634 199594 169662 199650
rect 169588 199566 169662 199594
rect 169484 196580 169536 196586
rect 169484 196522 169536 196528
rect 169588 196246 169616 199566
rect 169668 199504 169720 199510
rect 169668 199446 169720 199452
rect 169680 196489 169708 199446
rect 169772 197198 169800 199702
rect 169944 199718 169996 199724
rect 170128 199776 170180 199782
rect 170278 199764 170306 200124
rect 170128 199718 170180 199724
rect 170232 199736 170306 199764
rect 170370 199764 170398 200124
rect 170462 199918 170490 200124
rect 170554 199918 170582 200124
rect 170646 199923 170674 200124
rect 170450 199912 170502 199918
rect 170450 199854 170502 199860
rect 170542 199912 170594 199918
rect 170542 199854 170594 199860
rect 170632 199914 170688 199923
rect 170632 199849 170688 199858
rect 170496 199776 170548 199782
rect 170370 199736 170444 199764
rect 169850 199679 169906 199688
rect 169864 198626 169892 199679
rect 169852 198620 169904 198626
rect 169852 198562 169904 198568
rect 169760 197192 169812 197198
rect 169760 197134 169812 197140
rect 169760 196648 169812 196654
rect 169760 196590 169812 196596
rect 169666 196480 169722 196489
rect 169666 196415 169722 196424
rect 169576 196240 169628 196246
rect 169576 196182 169628 196188
rect 169668 195424 169720 195430
rect 169668 195366 169720 195372
rect 169680 195090 169708 195366
rect 169668 195084 169720 195090
rect 169668 195026 169720 195032
rect 169392 190256 169444 190262
rect 169392 190198 169444 190204
rect 169300 189644 169352 189650
rect 169300 189586 169352 189592
rect 169208 185768 169260 185774
rect 169208 185710 169260 185716
rect 168760 184742 168880 184770
rect 168760 184618 168788 184742
rect 168748 184612 168800 184618
rect 168748 184554 168800 184560
rect 168760 184006 168788 184554
rect 168748 184000 168800 184006
rect 168748 183942 168800 183948
rect 168656 180124 168708 180130
rect 168656 180066 168708 180072
rect 168564 148572 168616 148578
rect 168564 148514 168616 148520
rect 168470 148472 168526 148481
rect 168470 148407 168526 148416
rect 168380 147008 168432 147014
rect 168380 146950 168432 146956
rect 169772 146962 169800 196590
rect 169864 148510 169892 198562
rect 169956 195294 169984 199718
rect 170036 199708 170088 199714
rect 170036 199650 170088 199656
rect 170048 196654 170076 199650
rect 170036 196648 170088 196654
rect 170036 196590 170088 196596
rect 170140 196586 170168 199718
rect 170128 196580 170180 196586
rect 170128 196522 170180 196528
rect 169944 195288 169996 195294
rect 169944 195230 169996 195236
rect 169944 195016 169996 195022
rect 170232 194993 170260 199736
rect 170310 199608 170366 199617
rect 170310 199543 170366 199552
rect 170324 199374 170352 199543
rect 170312 199368 170364 199374
rect 170312 199310 170364 199316
rect 170312 196920 170364 196926
rect 170312 196862 170364 196868
rect 169944 194958 169996 194964
rect 170218 194984 170274 194993
rect 169956 184686 169984 194958
rect 170218 194919 170274 194928
rect 170324 189718 170352 196862
rect 170416 194274 170444 199736
rect 170496 199718 170548 199724
rect 170588 199776 170640 199782
rect 170738 199764 170766 200124
rect 170588 199718 170640 199724
rect 170692 199736 170766 199764
rect 170830 199764 170858 200124
rect 170922 199923 170950 200124
rect 170908 199914 170964 199923
rect 171014 199918 171042 200124
rect 170908 199849 170964 199858
rect 171002 199912 171054 199918
rect 171002 199854 171054 199860
rect 170956 199776 171008 199782
rect 170830 199736 170904 199764
rect 170508 196654 170536 199718
rect 170600 198422 170628 199718
rect 170588 198416 170640 198422
rect 170588 198358 170640 198364
rect 170588 197668 170640 197674
rect 170588 197610 170640 197616
rect 170496 196648 170548 196654
rect 170496 196590 170548 196596
rect 170496 195560 170548 195566
rect 170496 195502 170548 195508
rect 170404 194268 170456 194274
rect 170404 194210 170456 194216
rect 170508 193254 170536 195502
rect 170496 193248 170548 193254
rect 170496 193190 170548 193196
rect 170508 190330 170536 193190
rect 170496 190324 170548 190330
rect 170496 190266 170548 190272
rect 170312 189712 170364 189718
rect 170312 189654 170364 189660
rect 170034 187640 170090 187649
rect 170034 187575 170090 187584
rect 169944 184680 169996 184686
rect 169944 184622 169996 184628
rect 170048 184550 170076 187575
rect 170404 185836 170456 185842
rect 170404 185778 170456 185784
rect 170036 184544 170088 184550
rect 170036 184486 170088 184492
rect 170416 178906 170444 185778
rect 170404 178900 170456 178906
rect 170404 178842 170456 178848
rect 169852 148504 169904 148510
rect 169852 148446 169904 148452
rect 169772 146934 169984 146962
rect 169852 145920 169904 145926
rect 169852 145862 169904 145868
rect 167368 145852 167420 145858
rect 167368 145794 167420 145800
rect 166908 144764 166960 144770
rect 166908 144706 166960 144712
rect 166448 142860 166500 142866
rect 166448 142802 166500 142808
rect 165618 141808 165674 141817
rect 165618 141743 165674 141752
rect 165160 141568 165212 141574
rect 165160 141510 165212 141516
rect 164976 140752 165028 140758
rect 164976 140694 165028 140700
rect 164988 139890 165016 140694
rect 166460 139890 166488 142802
rect 164436 139862 164496 139890
rect 164988 139862 165324 139890
rect 166152 139862 166488 139890
rect 166920 139890 166948 144706
rect 167380 139890 167408 145794
rect 169022 145752 169078 145761
rect 169022 145687 169078 145696
rect 168932 142928 168984 142934
rect 168932 142870 168984 142876
rect 168944 139890 168972 142870
rect 166920 139862 166980 139890
rect 167380 139862 167808 139890
rect 168636 139862 168972 139890
rect 169036 139890 169064 145687
rect 169758 143576 169814 143585
rect 169758 143511 169814 143520
rect 169772 142866 169800 143511
rect 169760 142860 169812 142866
rect 169760 142802 169812 142808
rect 169864 139890 169892 145862
rect 169956 140214 169984 146934
rect 169944 140208 169996 140214
rect 169944 140150 169996 140156
rect 169036 139862 169464 139890
rect 169864 139862 170292 139890
rect 141606 139360 141662 139369
rect 128450 139295 128506 139304
rect 129004 139324 129056 139330
rect 141436 139318 141606 139346
rect 141606 139295 141662 139304
rect 146666 139360 146722 139369
rect 146666 139295 146722 139304
rect 154026 139360 154082 139369
rect 170600 139330 170628 197610
rect 170692 195022 170720 199736
rect 170876 199617 170904 199736
rect 171106 199764 171134 200124
rect 170956 199718 171008 199724
rect 171060 199736 171134 199764
rect 170862 199608 170918 199617
rect 170862 199543 170918 199552
rect 170772 199436 170824 199442
rect 170968 199424 170996 199718
rect 170772 199378 170824 199384
rect 170876 199396 170996 199424
rect 170784 197606 170812 199378
rect 170772 197600 170824 197606
rect 170876 197577 170904 199396
rect 170954 199336 171010 199345
rect 170954 199271 171010 199280
rect 170968 198801 170996 199271
rect 170954 198792 171010 198801
rect 170954 198727 171010 198736
rect 170772 197542 170824 197548
rect 170862 197568 170918 197577
rect 170862 197503 170918 197512
rect 170770 197432 170826 197441
rect 170770 197367 170826 197376
rect 170784 197266 170812 197367
rect 170864 197328 170916 197334
rect 170864 197270 170916 197276
rect 170772 197260 170824 197266
rect 170772 197202 170824 197208
rect 170876 196926 170904 197270
rect 170864 196920 170916 196926
rect 170770 196888 170826 196897
rect 170864 196862 170916 196868
rect 170770 196823 170772 196832
rect 170824 196823 170826 196832
rect 170772 196794 170824 196800
rect 170862 196752 170918 196761
rect 171060 196738 171088 199736
rect 171198 199696 171226 200124
rect 171290 199918 171318 200124
rect 171382 199918 171410 200124
rect 171474 199918 171502 200124
rect 171278 199912 171330 199918
rect 171278 199854 171330 199860
rect 171370 199912 171422 199918
rect 171370 199854 171422 199860
rect 171462 199912 171514 199918
rect 171462 199854 171514 199860
rect 171416 199776 171468 199782
rect 170862 196687 170918 196696
rect 170968 196710 171088 196738
rect 171152 199668 171226 199696
rect 171322 199744 171378 199753
rect 171566 199730 171594 200124
rect 171658 199923 171686 200124
rect 171644 199914 171700 199923
rect 171644 199849 171700 199858
rect 171416 199718 171468 199724
rect 171322 199679 171378 199688
rect 170876 195770 170904 196687
rect 170864 195764 170916 195770
rect 170864 195706 170916 195712
rect 170772 195696 170824 195702
rect 170968 195673 170996 196710
rect 171152 196636 171180 199668
rect 171232 199504 171284 199510
rect 171232 199446 171284 199452
rect 171060 196608 171180 196636
rect 170772 195638 170824 195644
rect 170954 195664 171010 195673
rect 170680 195016 170732 195022
rect 170680 194958 170732 194964
rect 170784 189582 170812 195638
rect 170954 195599 171010 195608
rect 170772 189576 170824 189582
rect 170772 189518 170824 189524
rect 171060 188562 171088 196608
rect 171140 196444 171192 196450
rect 171140 196386 171192 196392
rect 171048 188556 171100 188562
rect 171048 188498 171100 188504
rect 171152 161430 171180 196386
rect 171244 181966 171272 199446
rect 171336 195906 171364 199679
rect 171428 197674 171456 199718
rect 171520 199702 171594 199730
rect 171520 198558 171548 199702
rect 171750 199696 171778 200124
rect 171842 199918 171870 200124
rect 171934 199918 171962 200124
rect 172026 199923 172054 200124
rect 171830 199912 171882 199918
rect 171830 199854 171882 199860
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 172012 199914 172068 199923
rect 172012 199849 172068 199858
rect 171968 199776 172020 199782
rect 172118 199764 172146 200124
rect 172210 199782 172238 200124
rect 171968 199718 172020 199724
rect 172072 199736 172146 199764
rect 172198 199776 172250 199782
rect 171750 199668 171824 199696
rect 171690 199608 171746 199617
rect 171600 199572 171652 199578
rect 171690 199543 171746 199552
rect 171600 199514 171652 199520
rect 171508 198552 171560 198558
rect 171508 198494 171560 198500
rect 171416 197668 171468 197674
rect 171416 197610 171468 197616
rect 171508 197396 171560 197402
rect 171508 197338 171560 197344
rect 171416 197192 171468 197198
rect 171416 197134 171468 197140
rect 171324 195900 171376 195906
rect 171324 195842 171376 195848
rect 171428 194857 171456 197134
rect 171414 194848 171470 194857
rect 171414 194783 171470 194792
rect 171520 193798 171548 197338
rect 171612 197198 171640 199514
rect 171704 199073 171732 199543
rect 171796 199510 171824 199668
rect 171784 199504 171836 199510
rect 171980 199492 172008 199718
rect 171784 199446 171836 199452
rect 171888 199464 172008 199492
rect 171690 199064 171746 199073
rect 171690 198999 171746 199008
rect 171888 198812 171916 199464
rect 172072 199424 172100 199736
rect 172302 199764 172330 200124
rect 172394 199918 172422 200124
rect 172486 199923 172514 200124
rect 172382 199912 172434 199918
rect 172382 199854 172434 199860
rect 172472 199914 172528 199923
rect 172578 199918 172606 200124
rect 172472 199849 172528 199858
rect 172566 199912 172618 199918
rect 172566 199854 172618 199860
rect 172670 199764 172698 200124
rect 172762 199889 172790 200124
rect 172854 199918 172882 200124
rect 172946 199918 172974 200124
rect 173038 199918 173066 200124
rect 172842 199912 172894 199918
rect 172748 199880 172804 199889
rect 172842 199854 172894 199860
rect 172934 199912 172986 199918
rect 172934 199854 172986 199860
rect 173026 199912 173078 199918
rect 173130 199889 173158 200124
rect 173222 199918 173250 200124
rect 173210 199912 173262 199918
rect 173026 199854 173078 199860
rect 173116 199880 173172 199889
rect 172748 199815 172804 199824
rect 173210 199854 173262 199860
rect 173116 199815 173172 199824
rect 172796 199776 172848 199782
rect 172302 199736 172376 199764
rect 172670 199736 172744 199764
rect 172198 199718 172250 199724
rect 172152 199640 172204 199646
rect 172152 199582 172204 199588
rect 171796 198784 171916 198812
rect 171980 199396 172100 199424
rect 171796 198218 171824 198784
rect 171980 198734 172008 199396
rect 172164 199322 172192 199582
rect 172244 199572 172296 199578
rect 172244 199514 172296 199520
rect 171888 198706 172008 198734
rect 172072 199294 172192 199322
rect 171784 198212 171836 198218
rect 171784 198154 171836 198160
rect 171600 197192 171652 197198
rect 171888 197146 171916 198706
rect 171968 197260 172020 197266
rect 171968 197202 172020 197208
rect 171600 197134 171652 197140
rect 171704 197118 171916 197146
rect 171508 193792 171560 193798
rect 171508 193734 171560 193740
rect 171704 192642 171732 197118
rect 171980 196994 172008 197202
rect 171876 196988 171928 196994
rect 171876 196930 171928 196936
rect 171968 196988 172020 196994
rect 171968 196930 172020 196936
rect 171888 195106 171916 196930
rect 171968 196580 172020 196586
rect 171968 196522 172020 196528
rect 171796 195078 171916 195106
rect 171692 192636 171744 192642
rect 171692 192578 171744 192584
rect 171796 190330 171824 195078
rect 171876 194812 171928 194818
rect 171876 194754 171928 194760
rect 171784 190324 171836 190330
rect 171784 190266 171836 190272
rect 171232 181960 171284 181966
rect 171232 181902 171284 181908
rect 171140 161424 171192 161430
rect 171140 161366 171192 161372
rect 171888 147354 171916 194754
rect 171980 187678 172008 196522
rect 172072 196450 172100 199294
rect 172256 198150 172284 199514
rect 172348 198937 172376 199736
rect 172428 199708 172480 199714
rect 172428 199650 172480 199656
rect 172334 198928 172390 198937
rect 172334 198863 172390 198872
rect 172244 198144 172296 198150
rect 172244 198086 172296 198092
rect 172440 197962 172468 199650
rect 172612 199640 172664 199646
rect 172612 199582 172664 199588
rect 172624 199481 172652 199582
rect 172610 199472 172666 199481
rect 172610 199407 172666 199416
rect 172256 197934 172468 197962
rect 172060 196444 172112 196450
rect 172060 196386 172112 196392
rect 172256 192914 172284 197934
rect 172624 197826 172652 199407
rect 172440 197798 172652 197826
rect 172336 197260 172388 197266
rect 172336 197202 172388 197208
rect 172244 192908 172296 192914
rect 172244 192850 172296 192856
rect 171968 187672 172020 187678
rect 171968 187614 172020 187620
rect 172244 187672 172296 187678
rect 172244 187614 172296 187620
rect 172256 184618 172284 187614
rect 172244 184612 172296 184618
rect 172244 184554 172296 184560
rect 172244 161424 172296 161430
rect 172244 161366 172296 161372
rect 172256 160750 172284 161366
rect 172244 160744 172296 160750
rect 172244 160686 172296 160692
rect 172348 148238 172376 197202
rect 172336 148232 172388 148238
rect 172336 148174 172388 148180
rect 171876 147348 171928 147354
rect 171876 147290 171928 147296
rect 171506 145888 171562 145897
rect 171506 145823 171562 145832
rect 171048 142860 171100 142866
rect 171048 142802 171100 142808
rect 171060 139890 171088 142802
rect 171520 139890 171548 145823
rect 172440 141982 172468 197798
rect 172520 197736 172572 197742
rect 172520 197678 172572 197684
rect 172532 193225 172560 197678
rect 172716 197402 172744 199736
rect 172796 199718 172848 199724
rect 173164 199776 173216 199782
rect 173314 199764 173342 200124
rect 173164 199718 173216 199724
rect 173268 199736 173342 199764
rect 172704 197396 172756 197402
rect 172704 197338 172756 197344
rect 172518 193216 172574 193225
rect 172518 193151 172574 193160
rect 172808 191834 172836 199718
rect 172888 199708 172940 199714
rect 172888 199650 172940 199656
rect 172900 197742 172928 199650
rect 172980 199640 173032 199646
rect 172980 199582 173032 199588
rect 172992 198694 173020 199582
rect 172980 198688 173032 198694
rect 172980 198630 173032 198636
rect 173072 198552 173124 198558
rect 173072 198494 173124 198500
rect 172980 198212 173032 198218
rect 172980 198154 173032 198160
rect 172888 197736 172940 197742
rect 172888 197678 172940 197684
rect 172992 196489 173020 198154
rect 173084 196761 173112 198494
rect 173070 196752 173126 196761
rect 173070 196687 173126 196696
rect 172978 196480 173034 196489
rect 173176 196432 173204 199718
rect 173268 198665 173296 199736
rect 173406 199492 173434 200124
rect 173498 199918 173526 200124
rect 173486 199912 173538 199918
rect 173486 199854 173538 199860
rect 173590 199764 173618 200124
rect 173682 199918 173710 200124
rect 173670 199912 173722 199918
rect 173670 199854 173722 199860
rect 173774 199764 173802 200124
rect 173866 199923 173894 200124
rect 173852 199914 173908 199923
rect 173958 199918 173986 200124
rect 174050 199918 174078 200124
rect 174142 199918 174170 200124
rect 173852 199849 173908 199858
rect 173946 199912 173998 199918
rect 173946 199854 173998 199860
rect 174038 199912 174090 199918
rect 174038 199854 174090 199860
rect 174130 199912 174182 199918
rect 174130 199854 174182 199860
rect 173590 199736 173664 199764
rect 173532 199640 173584 199646
rect 173532 199582 173584 199588
rect 173360 199464 173434 199492
rect 173254 198656 173310 198665
rect 173254 198591 173310 198600
rect 173360 197266 173388 199464
rect 173440 198824 173492 198830
rect 173440 198766 173492 198772
rect 173348 197260 173400 197266
rect 173348 197202 173400 197208
rect 173346 197024 173402 197033
rect 173346 196959 173402 196968
rect 173360 196858 173388 196959
rect 173348 196852 173400 196858
rect 173348 196794 173400 196800
rect 173348 196648 173400 196654
rect 173348 196590 173400 196596
rect 172978 196415 173034 196424
rect 173084 196404 173204 196432
rect 172888 196376 172940 196382
rect 172888 196318 172940 196324
rect 172624 191806 172836 191834
rect 172624 191622 172652 191806
rect 172612 191616 172664 191622
rect 172612 191558 172664 191564
rect 172900 188290 172928 196318
rect 173084 195566 173112 196404
rect 173164 196308 173216 196314
rect 173164 196250 173216 196256
rect 173072 195560 173124 195566
rect 173072 195502 173124 195508
rect 172888 188284 172940 188290
rect 172888 188226 172940 188232
rect 172612 146056 172664 146062
rect 172612 145998 172664 146004
rect 172520 143540 172572 143546
rect 172520 143482 172572 143488
rect 172428 141976 172480 141982
rect 172428 141918 172480 141924
rect 172532 141438 172560 143482
rect 172520 141432 172572 141438
rect 172520 141374 172572 141380
rect 172624 139890 172652 145998
rect 173176 140350 173204 196250
rect 173256 192568 173308 192574
rect 173256 192510 173308 192516
rect 173268 142050 173296 192510
rect 173360 184754 173388 196590
rect 173452 195809 173480 198766
rect 173438 195800 173494 195809
rect 173438 195735 173494 195744
rect 173452 187134 173480 195735
rect 173544 195684 173572 199582
rect 173636 198830 173664 199736
rect 173728 199736 173802 199764
rect 173992 199776 174044 199782
rect 173852 199744 173908 199753
rect 173624 198824 173676 198830
rect 173624 198766 173676 198772
rect 173728 198665 173756 199736
rect 174234 199764 174262 200124
rect 174326 199923 174354 200124
rect 174312 199914 174368 199923
rect 174418 199918 174446 200124
rect 174510 199923 174538 200124
rect 174312 199849 174368 199858
rect 174406 199912 174458 199918
rect 174406 199854 174458 199860
rect 174496 199914 174552 199923
rect 174602 199918 174630 200124
rect 174694 199923 174722 200124
rect 174496 199849 174552 199858
rect 174590 199912 174642 199918
rect 174590 199854 174642 199860
rect 174680 199914 174736 199923
rect 174786 199918 174814 200124
rect 174680 199849 174736 199858
rect 174774 199912 174826 199918
rect 174774 199854 174826 199860
rect 174452 199776 174504 199782
rect 174234 199736 174400 199764
rect 173992 199718 174044 199724
rect 173852 199679 173854 199688
rect 173906 199679 173908 199688
rect 173854 199650 173906 199656
rect 173714 198656 173770 198665
rect 173714 198591 173770 198600
rect 173900 198144 173952 198150
rect 173900 198086 173952 198092
rect 173912 197266 173940 198086
rect 173900 197260 173952 197266
rect 173900 197202 173952 197208
rect 174004 196296 174032 199718
rect 174268 199572 174320 199578
rect 174268 199514 174320 199520
rect 174084 198688 174136 198694
rect 174084 198630 174136 198636
rect 174096 196926 174124 198630
rect 174084 196920 174136 196926
rect 174084 196862 174136 196868
rect 174084 196648 174136 196654
rect 174084 196590 174136 196596
rect 173912 196268 174032 196296
rect 173912 196110 173940 196268
rect 174096 196194 174124 196590
rect 174004 196166 174124 196194
rect 173900 196104 173952 196110
rect 173900 196046 173952 196052
rect 173900 195764 173952 195770
rect 173900 195706 173952 195712
rect 173544 195656 173848 195684
rect 173532 195560 173584 195566
rect 173532 195502 173584 195508
rect 173544 190454 173572 195502
rect 173714 193216 173770 193225
rect 173714 193151 173770 193160
rect 173728 190777 173756 193151
rect 173714 190768 173770 190777
rect 173714 190703 173770 190712
rect 173544 190426 173756 190454
rect 173440 187128 173492 187134
rect 173440 187070 173492 187076
rect 173348 184748 173400 184754
rect 173348 184690 173400 184696
rect 173728 143546 173756 190426
rect 173820 185842 173848 195656
rect 173912 195022 173940 195706
rect 173900 195016 173952 195022
rect 173900 194958 173952 194964
rect 173808 185836 173860 185842
rect 173808 185778 173860 185784
rect 174004 149054 174032 196166
rect 174084 196104 174136 196110
rect 174084 196046 174136 196052
rect 174176 196104 174228 196110
rect 174176 196046 174228 196052
rect 174096 181422 174124 196046
rect 174188 189922 174216 196046
rect 174280 192778 174308 199514
rect 174372 196654 174400 199736
rect 174728 199776 174780 199782
rect 174452 199718 174504 199724
rect 174542 199744 174598 199753
rect 174360 196648 174412 196654
rect 174360 196590 174412 196596
rect 174464 195838 174492 199718
rect 174728 199718 174780 199724
rect 174542 199679 174598 199688
rect 174636 199708 174688 199714
rect 174556 196081 174584 199679
rect 174636 199650 174688 199656
rect 174648 198898 174676 199650
rect 174636 198892 174688 198898
rect 174636 198834 174688 198840
rect 174634 198656 174690 198665
rect 174634 198591 174690 198600
rect 174542 196072 174598 196081
rect 174542 196007 174598 196016
rect 174452 195832 174504 195838
rect 174452 195774 174504 195780
rect 174360 195696 174412 195702
rect 174360 195638 174412 195644
rect 174372 194954 174400 195638
rect 174648 195106 174676 198591
rect 174740 195809 174768 199718
rect 174878 199696 174906 200124
rect 174970 199918 174998 200124
rect 175062 199918 175090 200124
rect 175154 199918 175182 200124
rect 175246 199918 175274 200124
rect 174958 199912 175010 199918
rect 174958 199854 175010 199860
rect 175050 199912 175102 199918
rect 175050 199854 175102 199860
rect 175142 199912 175194 199918
rect 175142 199854 175194 199860
rect 175234 199912 175286 199918
rect 175234 199854 175286 199860
rect 175338 199782 175366 200124
rect 175430 199918 175458 200124
rect 175418 199912 175470 199918
rect 175418 199854 175470 199860
rect 175096 199776 175148 199782
rect 175326 199776 175378 199782
rect 175148 199724 175228 199730
rect 175096 199718 175228 199724
rect 175522 199730 175550 200124
rect 175326 199718 175378 199724
rect 175108 199702 175228 199718
rect 174832 199668 174906 199696
rect 174832 196110 174860 199668
rect 175096 199640 175148 199646
rect 175096 199582 175148 199588
rect 174912 199572 174964 199578
rect 174912 199514 174964 199520
rect 175004 199572 175056 199578
rect 175004 199514 175056 199520
rect 174820 196104 174872 196110
rect 174820 196046 174872 196052
rect 174726 195800 174782 195809
rect 174726 195735 174782 195744
rect 174648 195078 174768 195106
rect 174636 195016 174688 195022
rect 174636 194958 174688 194964
rect 174360 194948 174412 194954
rect 174360 194890 174412 194896
rect 174544 194064 174596 194070
rect 174544 194006 174596 194012
rect 174268 192772 174320 192778
rect 174268 192714 174320 192720
rect 174176 189916 174228 189922
rect 174176 189858 174228 189864
rect 174084 181416 174136 181422
rect 174084 181358 174136 181364
rect 173992 149048 174044 149054
rect 173992 148990 174044 148996
rect 173992 146124 174044 146130
rect 173992 146066 174044 146072
rect 173716 143540 173768 143546
rect 173716 143482 173768 143488
rect 173728 142798 173756 143482
rect 173716 142792 173768 142798
rect 173716 142734 173768 142740
rect 173716 142520 173768 142526
rect 173716 142462 173768 142468
rect 173256 142044 173308 142050
rect 173256 141986 173308 141992
rect 173164 140344 173216 140350
rect 173164 140286 173216 140292
rect 173728 139890 173756 142462
rect 171060 139862 171120 139890
rect 171520 139862 171948 139890
rect 172624 139862 172776 139890
rect 173604 139862 173756 139890
rect 174004 139890 174032 146066
rect 174556 141370 174584 194006
rect 174648 148374 174676 194958
rect 174740 192681 174768 195078
rect 174726 192672 174782 192681
rect 174726 192607 174782 192616
rect 174924 191834 174952 199514
rect 175016 195702 175044 199514
rect 175004 195696 175056 195702
rect 175004 195638 175056 195644
rect 175108 192574 175136 199582
rect 175096 192568 175148 192574
rect 175096 192510 175148 192516
rect 175200 192438 175228 199702
rect 175476 199702 175550 199730
rect 175372 199640 175424 199646
rect 175372 199582 175424 199588
rect 175384 194594 175412 199582
rect 175476 195362 175504 199702
rect 175614 199594 175642 200124
rect 175706 199918 175734 200124
rect 175798 199923 175826 200124
rect 175694 199912 175746 199918
rect 175694 199854 175746 199860
rect 175784 199914 175840 199923
rect 175784 199849 175840 199858
rect 175890 199850 175918 200124
rect 175878 199844 175930 199850
rect 175878 199786 175930 199792
rect 175740 199708 175792 199714
rect 175740 199650 175792 199656
rect 175832 199708 175884 199714
rect 175832 199650 175884 199656
rect 175614 199566 175688 199594
rect 175556 198960 175608 198966
rect 175556 198902 175608 198908
rect 175464 195356 175516 195362
rect 175464 195298 175516 195304
rect 175292 194566 175412 194594
rect 175188 192432 175240 192438
rect 175188 192374 175240 192380
rect 174924 191806 175044 191834
rect 175016 180794 175044 191806
rect 174832 180766 175044 180794
rect 174636 148368 174688 148374
rect 174636 148310 174688 148316
rect 174832 141438 174860 180766
rect 175292 144838 175320 194566
rect 175568 193214 175596 198902
rect 175660 198626 175688 199566
rect 175648 198620 175700 198626
rect 175648 198562 175700 198568
rect 175752 197441 175780 199650
rect 175844 198966 175872 199650
rect 175982 199628 176010 200124
rect 176074 199764 176102 200124
rect 176166 199918 176194 200124
rect 176154 199912 176206 199918
rect 176154 199854 176206 199860
rect 176258 199764 176286 200124
rect 176350 199850 176378 200124
rect 176338 199844 176390 199850
rect 176338 199786 176390 199792
rect 176074 199736 176148 199764
rect 175936 199600 176010 199628
rect 175832 198960 175884 198966
rect 175832 198902 175884 198908
rect 175738 197432 175794 197441
rect 175738 197367 175794 197376
rect 175384 193186 175596 193214
rect 175384 148442 175412 193186
rect 175462 189136 175518 189145
rect 175462 189071 175518 189080
rect 175476 181354 175504 189071
rect 175646 186144 175702 186153
rect 175646 186079 175702 186088
rect 175660 185026 175688 186079
rect 175648 185020 175700 185026
rect 175648 184962 175700 184968
rect 175464 181348 175516 181354
rect 175464 181290 175516 181296
rect 175936 180794 175964 199600
rect 176120 197418 176148 199736
rect 176212 199736 176286 199764
rect 176442 199764 176470 200124
rect 176534 199918 176562 200124
rect 176626 199923 176654 200124
rect 176522 199912 176574 199918
rect 176522 199854 176574 199860
rect 176612 199914 176668 199923
rect 176718 199918 176746 200124
rect 176612 199849 176668 199858
rect 176706 199912 176758 199918
rect 176706 199854 176758 199860
rect 176810 199764 176838 200124
rect 176902 199923 176930 200124
rect 176888 199914 176944 199923
rect 176888 199849 176944 199858
rect 176994 199764 177022 200124
rect 176442 199736 176516 199764
rect 176212 199481 176240 199736
rect 176292 199640 176344 199646
rect 176292 199582 176344 199588
rect 176384 199640 176436 199646
rect 176384 199582 176436 199588
rect 176198 199472 176254 199481
rect 176198 199407 176254 199416
rect 176200 198960 176252 198966
rect 176200 198902 176252 198908
rect 176028 197390 176148 197418
rect 176028 194206 176056 197390
rect 176212 196432 176240 198902
rect 176304 196450 176332 199582
rect 176120 196404 176240 196432
rect 176292 196444 176344 196450
rect 176016 194200 176068 194206
rect 176016 194142 176068 194148
rect 176120 191554 176148 196404
rect 176292 196386 176344 196392
rect 176200 196172 176252 196178
rect 176200 196114 176252 196120
rect 176108 191548 176160 191554
rect 176108 191490 176160 191496
rect 175476 180766 175964 180794
rect 175476 151298 175504 180766
rect 175464 151292 175516 151298
rect 175464 151234 175516 151240
rect 175372 148436 175424 148442
rect 175372 148378 175424 148384
rect 176212 147286 176240 196114
rect 176292 195832 176344 195838
rect 176292 195774 176344 195780
rect 176304 195430 176332 195774
rect 176292 195424 176344 195430
rect 176292 195366 176344 195372
rect 176396 193225 176424 199582
rect 176488 199050 176516 199736
rect 176764 199736 176838 199764
rect 176948 199736 177022 199764
rect 176660 199504 176712 199510
rect 176660 199446 176712 199452
rect 176488 199022 176608 199050
rect 176580 198966 176608 199022
rect 176568 198960 176620 198966
rect 176568 198902 176620 198908
rect 176382 193216 176438 193225
rect 176382 193151 176438 193160
rect 176566 178664 176622 178673
rect 176566 178599 176622 178608
rect 176200 147280 176252 147286
rect 176200 147222 176252 147228
rect 176580 146985 176608 178599
rect 176566 146976 176622 146985
rect 176566 146911 176622 146920
rect 176672 144906 176700 199446
rect 176764 190454 176792 199736
rect 176948 199510 176976 199736
rect 177086 199696 177114 200124
rect 177178 199918 177206 200124
rect 177166 199912 177218 199918
rect 177166 199854 177218 199860
rect 177040 199668 177114 199696
rect 176936 199504 176988 199510
rect 176936 199446 176988 199452
rect 177040 198558 177068 199668
rect 177270 199628 177298 200124
rect 177362 199918 177390 200124
rect 177350 199912 177402 199918
rect 177350 199854 177402 199860
rect 177454 199730 177482 200124
rect 177546 199866 177574 200124
rect 177868 200110 178356 200138
rect 178130 200016 178186 200025
rect 178130 199951 178186 199960
rect 177854 199880 177910 199889
rect 177546 199838 177620 199866
rect 177224 199600 177298 199628
rect 177408 199702 177482 199730
rect 177028 198552 177080 198558
rect 177028 198494 177080 198500
rect 177120 194336 177172 194342
rect 177120 194278 177172 194284
rect 177132 194070 177160 194278
rect 177120 194064 177172 194070
rect 177120 194006 177172 194012
rect 176764 190426 176884 190454
rect 176752 186924 176804 186930
rect 176752 186866 176804 186872
rect 176764 184074 176792 186866
rect 176752 184068 176804 184074
rect 176752 184010 176804 184016
rect 176856 181898 176884 190426
rect 177224 188630 177252 199600
rect 177408 197033 177436 199702
rect 177488 197940 177540 197946
rect 177488 197882 177540 197888
rect 177394 197024 177450 197033
rect 177394 196959 177450 196968
rect 177212 188624 177264 188630
rect 177212 188566 177264 188572
rect 176844 181892 176896 181898
rect 176844 181834 176896 181840
rect 177304 145512 177356 145518
rect 177304 145454 177356 145460
rect 176660 144900 176712 144906
rect 176660 144842 176712 144848
rect 175280 144832 175332 144838
rect 175280 144774 175332 144780
rect 177212 143268 177264 143274
rect 177212 143210 177264 143216
rect 175188 143200 175240 143206
rect 175188 143142 175240 143148
rect 174820 141432 174872 141438
rect 174820 141374 174872 141380
rect 174544 141364 174596 141370
rect 174544 141306 174596 141312
rect 175200 139890 175228 143142
rect 176384 142724 176436 142730
rect 176384 142666 176436 142672
rect 176396 139890 176424 142666
rect 177224 142390 177252 143210
rect 177212 142384 177264 142390
rect 177212 142326 177264 142332
rect 177224 139890 177252 142326
rect 174004 139862 174432 139890
rect 175200 139862 175260 139890
rect 176088 139862 176424 139890
rect 176916 139862 177252 139890
rect 177316 139890 177344 145454
rect 177500 144158 177528 197882
rect 177592 197810 177620 199838
rect 177854 199815 177910 199824
rect 178040 199844 178092 199850
rect 177672 199776 177724 199782
rect 177672 199718 177724 199724
rect 177684 198801 177712 199718
rect 177764 198892 177816 198898
rect 177764 198834 177816 198840
rect 177670 198792 177726 198801
rect 177670 198727 177726 198736
rect 177672 198416 177724 198422
rect 177672 198358 177724 198364
rect 177580 197804 177632 197810
rect 177580 197746 177632 197752
rect 177580 197668 177632 197674
rect 177580 197610 177632 197616
rect 177592 146198 177620 197610
rect 177684 186862 177712 198358
rect 177776 188494 177804 198834
rect 177868 194070 177896 199815
rect 178040 199786 178092 199792
rect 178052 198966 178080 199786
rect 178040 198960 178092 198966
rect 178040 198902 178092 198908
rect 178144 195498 178172 199951
rect 178224 197804 178276 197810
rect 178224 197746 178276 197752
rect 178132 195492 178184 195498
rect 178132 195434 178184 195440
rect 178040 195220 178092 195226
rect 178040 195162 178092 195168
rect 178052 194614 178080 195162
rect 178040 194608 178092 194614
rect 178040 194550 178092 194556
rect 177856 194064 177908 194070
rect 177856 194006 177908 194012
rect 178052 193474 178080 194550
rect 178052 193446 178172 193474
rect 178040 193384 178092 193390
rect 178040 193326 178092 193332
rect 177764 188488 177816 188494
rect 177764 188430 177816 188436
rect 177672 186856 177724 186862
rect 177672 186798 177724 186804
rect 177580 146192 177632 146198
rect 177580 146134 177632 146140
rect 177488 144152 177540 144158
rect 177488 144094 177540 144100
rect 178052 141681 178080 193326
rect 178038 141672 178094 141681
rect 178038 141607 178094 141616
rect 178144 141506 178172 193446
rect 178236 185586 178264 197746
rect 178328 185858 178356 200110
rect 178408 200116 178460 200122
rect 178408 200058 178460 200064
rect 178420 198218 178448 200058
rect 178590 199744 178646 199753
rect 178590 199679 178646 199688
rect 178408 198212 178460 198218
rect 178408 198154 178460 198160
rect 178408 196444 178460 196450
rect 178408 196386 178460 196392
rect 178420 185978 178448 196386
rect 178604 194177 178632 199679
rect 178696 198937 178724 200398
rect 178774 200359 178830 200368
rect 178788 200258 178816 200359
rect 180430 200288 180486 200297
rect 178776 200252 178828 200258
rect 180430 200223 180486 200232
rect 178776 200194 178828 200200
rect 180062 200016 180118 200025
rect 180062 199951 180118 199960
rect 178960 199640 179012 199646
rect 178866 199608 178922 199617
rect 178960 199582 179012 199588
rect 178866 199543 178922 199552
rect 178682 198928 178738 198937
rect 178682 198863 178738 198872
rect 178684 196512 178736 196518
rect 178684 196454 178736 196460
rect 178590 194168 178646 194177
rect 178590 194103 178646 194112
rect 178408 185972 178460 185978
rect 178408 185914 178460 185920
rect 178328 185830 178448 185858
rect 178236 185558 178356 185586
rect 178224 183524 178276 183530
rect 178224 183466 178276 183472
rect 178236 183326 178264 183466
rect 178328 183462 178356 185558
rect 178420 183530 178448 185830
rect 178408 183524 178460 183530
rect 178408 183466 178460 183472
rect 178316 183456 178368 183462
rect 178316 183398 178368 183404
rect 178224 183320 178276 183326
rect 178224 183262 178276 183268
rect 178328 183258 178356 183398
rect 178316 183252 178368 183258
rect 178316 183194 178368 183200
rect 178590 143440 178646 143449
rect 178590 143375 178646 143384
rect 178604 142730 178632 143375
rect 178592 142724 178644 142730
rect 178592 142666 178644 142672
rect 178132 141500 178184 141506
rect 178132 141442 178184 141448
rect 178696 140554 178724 196454
rect 178776 194880 178828 194886
rect 178776 194822 178828 194828
rect 178684 140548 178736 140554
rect 178684 140490 178736 140496
rect 178788 140418 178816 194822
rect 178880 193390 178908 199543
rect 178972 198830 179000 199582
rect 179326 199472 179382 199481
rect 179326 199407 179382 199416
rect 178960 198824 179012 198830
rect 178960 198766 179012 198772
rect 179340 195566 179368 199407
rect 179602 199064 179658 199073
rect 179602 198999 179658 199008
rect 179512 198824 179564 198830
rect 179512 198766 179564 198772
rect 179418 197976 179474 197985
rect 179418 197911 179474 197920
rect 179328 195560 179380 195566
rect 179328 195502 179380 195508
rect 178868 193384 178920 193390
rect 178868 193326 178920 193332
rect 179326 191040 179382 191049
rect 179326 190975 179382 190984
rect 179340 151814 179368 190975
rect 179432 188698 179460 197911
rect 179420 188692 179472 188698
rect 179420 188634 179472 188640
rect 179248 151786 179368 151814
rect 178866 142896 178922 142905
rect 178866 142831 178922 142840
rect 178776 140412 178828 140418
rect 178776 140354 178828 140360
rect 178880 139890 178908 142831
rect 179248 140321 179276 151786
rect 179328 143404 179380 143410
rect 179328 143346 179380 143352
rect 179234 140312 179290 140321
rect 179234 140247 179290 140256
rect 177316 139862 177744 139890
rect 178572 139862 178908 139890
rect 179340 139890 179368 143346
rect 179418 143032 179474 143041
rect 179418 142967 179474 142976
rect 179432 142526 179460 142967
rect 179420 142520 179472 142526
rect 179420 142462 179472 142468
rect 179524 141545 179552 198766
rect 179510 141536 179566 141545
rect 179510 141471 179566 141480
rect 179616 141409 179644 198999
rect 180076 198529 180104 199951
rect 180444 199918 180472 200223
rect 180522 200152 180578 200161
rect 180522 200087 180578 200096
rect 180536 200054 180564 200087
rect 180524 200048 180576 200054
rect 180524 199990 180576 199996
rect 181812 199980 181864 199986
rect 181812 199922 181864 199928
rect 180432 199912 180484 199918
rect 180432 199854 180484 199860
rect 180246 199744 180302 199753
rect 180246 199679 180302 199688
rect 180062 198520 180118 198529
rect 180062 198455 180118 198464
rect 179880 146260 179932 146266
rect 179880 146202 179932 146208
rect 179696 142792 179748 142798
rect 179696 142734 179748 142740
rect 179708 142526 179736 142734
rect 179696 142520 179748 142526
rect 179696 142462 179748 142468
rect 179602 141400 179658 141409
rect 179602 141335 179658 141344
rect 179892 139890 179920 146202
rect 180076 140486 180104 198455
rect 180260 198393 180288 199679
rect 180706 199472 180762 199481
rect 180706 199407 180762 199416
rect 180720 199073 180748 199407
rect 180706 199064 180762 199073
rect 180706 198999 180762 199008
rect 180246 198384 180302 198393
rect 180246 198319 180302 198328
rect 180156 195084 180208 195090
rect 180156 195026 180208 195032
rect 180168 140622 180196 195026
rect 180260 148170 180288 198319
rect 181824 195129 181852 199922
rect 188988 199776 189040 199782
rect 188988 199718 189040 199724
rect 182272 199708 182324 199714
rect 182272 199650 182324 199656
rect 182180 199368 182232 199374
rect 182180 199310 182232 199316
rect 182192 198150 182220 199310
rect 182284 198694 182312 199650
rect 184756 199572 184808 199578
rect 184756 199514 184808 199520
rect 182272 198688 182324 198694
rect 182272 198630 182324 198636
rect 183560 198484 183612 198490
rect 183560 198426 183612 198432
rect 182180 198144 182232 198150
rect 182180 198086 182232 198092
rect 183572 197985 183600 198426
rect 183558 197976 183614 197985
rect 183558 197911 183614 197920
rect 182824 195152 182876 195158
rect 181810 195120 181866 195129
rect 182824 195094 182876 195100
rect 181810 195055 181866 195064
rect 182086 191448 182142 191457
rect 182086 191383 182142 191392
rect 182100 191185 182128 191383
rect 182086 191176 182142 191185
rect 182086 191111 182142 191120
rect 181996 187060 182048 187066
rect 181996 187002 182048 187008
rect 181904 184272 181956 184278
rect 181904 184214 181956 184220
rect 180708 181688 180760 181694
rect 180708 181630 180760 181636
rect 180616 178696 180668 178702
rect 180616 178638 180668 178644
rect 180248 148164 180300 148170
rect 180248 148106 180300 148112
rect 180628 142154 180656 178638
rect 180536 142126 180656 142154
rect 180156 140616 180208 140622
rect 180156 140558 180208 140564
rect 180064 140480 180116 140486
rect 180064 140422 180116 140428
rect 179340 139862 179400 139890
rect 179892 139862 180228 139890
rect 180536 139369 180564 142126
rect 180720 139369 180748 181630
rect 181444 145444 181496 145450
rect 181444 145386 181496 145392
rect 181352 143336 181404 143342
rect 181352 143278 181404 143284
rect 181364 139890 181392 143278
rect 181056 139862 181392 139890
rect 181456 139890 181484 145386
rect 181916 141681 181944 184214
rect 182008 141953 182036 187002
rect 181994 141944 182050 141953
rect 181994 141879 182050 141888
rect 181902 141672 181958 141681
rect 181902 141607 181958 141616
rect 181456 139862 181884 139890
rect 182100 139482 182128 191111
rect 182270 146024 182326 146033
rect 182270 145959 182326 145968
rect 182284 139890 182312 145959
rect 182836 140758 182864 195094
rect 183468 191140 183520 191146
rect 183468 191082 183520 191088
rect 183374 184512 183430 184521
rect 183374 184447 183430 184456
rect 183284 146872 183336 146878
rect 183284 146814 183336 146820
rect 182824 140752 182876 140758
rect 182824 140694 182876 140700
rect 183296 140593 183324 146814
rect 183388 141545 183416 184447
rect 183480 146878 183508 191082
rect 183468 146872 183520 146878
rect 183468 146814 183520 146820
rect 184768 144401 184796 199514
rect 184940 199504 184992 199510
rect 184940 199446 184992 199452
rect 186228 199504 186280 199510
rect 186228 199446 186280 199452
rect 184952 199102 184980 199446
rect 184940 199096 184992 199102
rect 184940 199038 184992 199044
rect 185400 198892 185452 198898
rect 185400 198834 185452 198840
rect 184848 198756 184900 198762
rect 184848 198698 184900 198704
rect 184754 144392 184810 144401
rect 184754 144327 184810 144336
rect 183466 142760 183522 142769
rect 183466 142695 183522 142704
rect 183374 141536 183430 141545
rect 183374 141471 183430 141480
rect 183282 140584 183338 140593
rect 183282 140519 183338 140528
rect 183480 139890 183508 142695
rect 184662 142624 184718 142633
rect 184662 142559 184718 142568
rect 184676 139890 184704 142559
rect 184860 140729 184888 198698
rect 185412 196654 185440 198834
rect 185400 196648 185452 196654
rect 185400 196590 185452 196596
rect 185584 193724 185636 193730
rect 185584 193666 185636 193672
rect 184940 145376 184992 145382
rect 184940 145318 184992 145324
rect 184846 140720 184902 140729
rect 184846 140655 184902 140664
rect 182284 139862 182712 139890
rect 183480 139862 183540 139890
rect 184368 139862 184704 139890
rect 184952 139890 184980 145318
rect 185596 140010 185624 193666
rect 185676 191480 185728 191486
rect 185676 191422 185728 191428
rect 185688 173194 185716 191422
rect 186136 189780 186188 189786
rect 186136 189722 186188 189728
rect 185676 173188 185728 173194
rect 185676 173130 185728 173136
rect 185688 171134 185716 173130
rect 185688 171106 186084 171134
rect 186056 151814 186084 171106
rect 185872 151786 186084 151814
rect 185584 140004 185636 140010
rect 185584 139946 185636 139952
rect 185872 139942 185900 151786
rect 186148 147098 186176 189722
rect 185964 147070 186176 147098
rect 185964 140690 185992 147070
rect 186240 146962 186268 199446
rect 188620 193792 188672 193798
rect 188620 193734 188672 193740
rect 186412 191412 186464 191418
rect 186412 191354 186464 191360
rect 186148 146934 186268 146962
rect 185952 140684 186004 140690
rect 185952 140626 186004 140632
rect 186148 140457 186176 146934
rect 186226 143168 186282 143177
rect 186226 143103 186282 143112
rect 186134 140448 186190 140457
rect 186134 140383 186190 140392
rect 185860 139936 185912 139942
rect 184952 139862 185196 139890
rect 186240 139890 186268 143103
rect 186320 140276 186372 140282
rect 186320 140218 186372 140224
rect 185860 139878 185912 139884
rect 186024 139862 186268 139890
rect 186332 139505 186360 140218
rect 182178 139496 182234 139505
rect 182100 139454 182178 139482
rect 182178 139431 182234 139440
rect 186318 139496 186374 139505
rect 186318 139431 186374 139440
rect 186424 139369 186452 191354
rect 187146 191176 187202 191185
rect 187146 191111 187202 191120
rect 187160 190913 187188 191111
rect 187146 190904 187202 190913
rect 187146 190839 187202 190848
rect 187056 188420 187108 188426
rect 187056 188362 187108 188368
rect 186778 143440 186834 143449
rect 186778 143375 186834 143384
rect 186962 143440 187018 143449
rect 186962 143375 187018 143384
rect 186792 143041 186820 143375
rect 186594 143032 186650 143041
rect 186594 142967 186650 142976
rect 186778 143032 186834 143041
rect 186778 142967 186834 142976
rect 186608 142497 186636 142967
rect 186594 142488 186650 142497
rect 186594 142423 186650 142432
rect 186976 139890 187004 143375
rect 186852 139862 187004 139890
rect 187068 139369 187096 188362
rect 187160 139777 187188 190839
rect 187516 182232 187568 182238
rect 187516 182174 187568 182180
rect 187528 147674 187556 182174
rect 188344 164280 188396 164286
rect 188344 164222 188396 164228
rect 188356 151814 188384 164222
rect 187436 147646 187556 147674
rect 188172 151786 188384 151814
rect 187146 139768 187202 139777
rect 187146 139703 187202 139712
rect 187436 139641 187464 147646
rect 187514 144256 187570 144265
rect 188172 144226 188200 151786
rect 188344 145988 188396 145994
rect 188344 145930 188396 145936
rect 188252 145036 188304 145042
rect 188252 144978 188304 144984
rect 187514 144191 187570 144200
rect 188160 144220 188212 144226
rect 187422 139632 187478 139641
rect 187422 139567 187478 139576
rect 187528 139505 187556 144191
rect 188160 144162 188212 144168
rect 187608 144084 187660 144090
rect 187608 144026 187660 144032
rect 187620 143410 187648 144026
rect 187608 143404 187660 143410
rect 187608 143346 187660 143352
rect 187606 143168 187662 143177
rect 187606 143103 187662 143112
rect 187620 142390 187648 143103
rect 187608 142384 187660 142390
rect 187608 142326 187660 142332
rect 187620 139890 187648 142326
rect 187620 139862 187680 139890
rect 187514 139496 187570 139505
rect 187514 139431 187570 139440
rect 180522 139360 180578 139369
rect 154026 139295 154082 139304
rect 170588 139324 170640 139330
rect 129004 139266 129056 139272
rect 180522 139295 180578 139304
rect 180706 139360 180762 139369
rect 180706 139295 180762 139304
rect 186410 139360 186466 139369
rect 186410 139295 186466 139304
rect 187054 139360 187110 139369
rect 188264 139330 188292 144978
rect 188356 139874 188384 145930
rect 188344 139868 188396 139874
rect 188344 139810 188396 139816
rect 187054 139295 187110 139304
rect 188252 139324 188304 139330
rect 170588 139266 170640 139272
rect 188252 139266 188304 139272
rect 188632 81734 188660 193734
rect 188712 193248 188764 193254
rect 188712 193190 188764 193196
rect 188620 81728 188672 81734
rect 188620 81670 188672 81676
rect 188620 81048 188672 81054
rect 188620 80990 188672 80996
rect 131764 80708 131816 80714
rect 131764 80650 131816 80656
rect 131856 80708 131908 80714
rect 132040 80708 132092 80714
rect 131908 80668 132040 80696
rect 131856 80650 131908 80656
rect 132040 80650 132092 80656
rect 177856 80708 177908 80714
rect 177856 80650 177908 80656
rect 177948 80708 178000 80714
rect 177948 80650 178000 80656
rect 182824 80708 182876 80714
rect 182824 80650 182876 80656
rect 123482 80608 123538 80617
rect 123482 80543 123538 80552
rect 122840 79620 122892 79626
rect 122840 79562 122892 79568
rect 122286 78568 122342 78577
rect 122286 78503 122342 78512
rect 122300 78266 122328 78503
rect 122288 78260 122340 78266
rect 122288 78202 122340 78208
rect 122852 68814 122880 79562
rect 123496 71777 123524 80543
rect 131776 80510 131804 80650
rect 123576 80504 123628 80510
rect 123576 80446 123628 80452
rect 131764 80504 131816 80510
rect 131764 80446 131816 80452
rect 123588 73166 123616 80446
rect 126244 80436 126296 80442
rect 126244 80378 126296 80384
rect 124588 80028 124640 80034
rect 124588 79970 124640 79976
rect 124600 78441 124628 79970
rect 125232 79892 125284 79898
rect 125232 79834 125284 79840
rect 124586 78432 124642 78441
rect 124586 78367 124642 78376
rect 125244 78130 125272 79834
rect 125232 78124 125284 78130
rect 125232 78066 125284 78072
rect 123576 73160 123628 73166
rect 123576 73102 123628 73108
rect 123482 71768 123538 71777
rect 123482 71703 123538 71712
rect 126256 71534 126284 80378
rect 126336 80368 126388 80374
rect 126336 80310 126388 80316
rect 128452 80368 128504 80374
rect 131856 80368 131908 80374
rect 128452 80310 128504 80316
rect 131854 80336 131856 80345
rect 131908 80336 131910 80345
rect 126348 72962 126376 80310
rect 127438 79792 127494 79801
rect 127438 79727 127494 79736
rect 127452 78538 127480 79727
rect 127532 79552 127584 79558
rect 127532 79494 127584 79500
rect 127440 78532 127492 78538
rect 127440 78474 127492 78480
rect 127544 74458 127572 79494
rect 128464 78577 128492 80310
rect 128636 80300 128688 80306
rect 131854 80271 131910 80280
rect 128636 80242 128688 80248
rect 128544 80232 128596 80238
rect 128544 80174 128596 80180
rect 128450 78568 128506 78577
rect 128450 78503 128506 78512
rect 128556 78402 128584 80174
rect 128544 78396 128596 78402
rect 128544 78338 128596 78344
rect 128648 78305 128676 80242
rect 132224 80232 132276 80238
rect 132222 80200 132224 80209
rect 177764 80232 177816 80238
rect 132276 80200 132278 80209
rect 132040 80164 132092 80170
rect 177764 80174 177816 80180
rect 132222 80135 132278 80144
rect 132040 80106 132092 80112
rect 131854 80064 131910 80073
rect 131854 79999 131910 80008
rect 129004 79688 129056 79694
rect 129002 79656 129004 79665
rect 129056 79656 129058 79665
rect 129002 79591 129058 79600
rect 131304 79620 131356 79626
rect 131304 79562 131356 79568
rect 129280 79484 129332 79490
rect 129280 79426 129332 79432
rect 128634 78296 128690 78305
rect 128634 78231 128690 78240
rect 128452 78056 128504 78062
rect 128452 77998 128504 78004
rect 129004 78056 129056 78062
rect 129004 77998 129056 78004
rect 128464 74497 128492 77998
rect 128450 74488 128506 74497
rect 127532 74452 127584 74458
rect 128450 74423 128506 74432
rect 127532 74394 127584 74400
rect 126336 72956 126388 72962
rect 126336 72898 126388 72904
rect 126244 71528 126296 71534
rect 126244 71470 126296 71476
rect 125600 70440 125652 70446
rect 125600 70382 125652 70388
rect 122196 68808 122248 68814
rect 122196 68750 122248 68756
rect 122840 68808 122892 68814
rect 122840 68750 122892 68756
rect 122104 64388 122156 64394
rect 122104 64330 122156 64336
rect 122208 41410 122236 68750
rect 122196 41404 122248 41410
rect 122196 41346 122248 41352
rect 117332 16546 117912 16574
rect 116584 4820 116636 4826
rect 116584 4762 116636 4768
rect 117884 480 117912 16546
rect 125612 480 125640 70382
rect 129016 65550 129044 77998
rect 129292 73166 129320 79426
rect 129648 78736 129700 78742
rect 129648 78678 129700 78684
rect 129660 78470 129688 78678
rect 131028 78600 131080 78606
rect 131028 78542 131080 78548
rect 129648 78464 129700 78470
rect 129648 78406 129700 78412
rect 129648 76628 129700 76634
rect 129648 76570 129700 76576
rect 129660 75818 129688 76570
rect 130384 75948 130436 75954
rect 130384 75890 130436 75896
rect 129648 75812 129700 75818
rect 129648 75754 129700 75760
rect 129280 73160 129332 73166
rect 129280 73102 129332 73108
rect 128452 65544 128504 65550
rect 128452 65486 128504 65492
rect 129004 65544 129056 65550
rect 129004 65486 129056 65492
rect 128360 64320 128412 64326
rect 128360 64262 128412 64268
rect 128372 16574 128400 64262
rect 128464 37262 128492 65486
rect 128452 37256 128504 37262
rect 128452 37198 128504 37204
rect 128372 16546 129504 16574
rect 129476 480 129504 16546
rect 130396 12442 130424 75890
rect 131040 72729 131068 78542
rect 131120 78464 131172 78470
rect 131120 78406 131172 78412
rect 131026 72720 131082 72729
rect 131026 72655 131082 72664
rect 131132 69018 131160 78406
rect 131212 78396 131264 78402
rect 131212 78338 131264 78344
rect 131224 73574 131252 78338
rect 131316 78334 131344 79562
rect 131868 78538 131896 79999
rect 131856 78532 131908 78538
rect 131856 78474 131908 78480
rect 131304 78328 131356 78334
rect 131304 78270 131356 78276
rect 132052 73778 132080 80106
rect 132328 80022 132388 80050
rect 132328 78470 132356 80022
rect 132466 79744 132494 80036
rect 132558 79966 132586 80036
rect 132650 79971 132678 80036
rect 132546 79960 132598 79966
rect 132546 79902 132598 79908
rect 132636 79962 132692 79971
rect 132636 79897 132692 79906
rect 132420 79716 132494 79744
rect 132592 79756 132644 79762
rect 132316 78464 132368 78470
rect 132316 78406 132368 78412
rect 132316 78124 132368 78130
rect 132316 78066 132368 78072
rect 132132 77308 132184 77314
rect 132132 77250 132184 77256
rect 132144 75070 132172 77250
rect 132132 75064 132184 75070
rect 132132 75006 132184 75012
rect 132040 73772 132092 73778
rect 132040 73714 132092 73720
rect 131212 73568 131264 73574
rect 131212 73510 131264 73516
rect 132328 73098 132356 78066
rect 132420 74526 132448 79716
rect 132592 79698 132644 79704
rect 132498 79656 132554 79665
rect 132498 79591 132554 79600
rect 132512 78470 132540 79591
rect 132500 78464 132552 78470
rect 132500 78406 132552 78412
rect 132604 75993 132632 79698
rect 132742 79676 132770 80036
rect 132834 79801 132862 80036
rect 132926 79966 132954 80036
rect 133018 79966 133046 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 132820 79792 132876 79801
rect 133110 79778 133138 80036
rect 133202 79971 133230 80036
rect 133188 79962 133244 79971
rect 133188 79897 133244 79906
rect 133294 79830 133322 80036
rect 133386 79966 133414 80036
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 132820 79727 132876 79736
rect 132972 79750 133138 79778
rect 133282 79824 133334 79830
rect 133478 79812 133506 80036
rect 133570 79830 133598 80036
rect 133662 79830 133690 80036
rect 133282 79766 133334 79772
rect 133432 79784 133506 79812
rect 133558 79824 133610 79830
rect 132742 79648 132816 79676
rect 132684 76152 132736 76158
rect 132684 76094 132736 76100
rect 132590 75984 132646 75993
rect 132590 75919 132646 75928
rect 132408 74520 132460 74526
rect 132408 74462 132460 74468
rect 131212 73092 131264 73098
rect 131212 73034 131264 73040
rect 132316 73092 132368 73098
rect 132316 73034 132368 73040
rect 131120 69012 131172 69018
rect 131120 68954 131172 68960
rect 131224 16590 131252 73034
rect 132696 67289 132724 76094
rect 132788 69562 132816 79648
rect 132866 79656 132922 79665
rect 132866 79591 132922 79600
rect 132880 76158 132908 79591
rect 132868 76152 132920 76158
rect 132868 76094 132920 76100
rect 132868 76016 132920 76022
rect 132868 75958 132920 75964
rect 132776 69556 132828 69562
rect 132776 69498 132828 69504
rect 132682 67280 132738 67289
rect 132682 67215 132738 67224
rect 132500 65408 132552 65414
rect 132500 65350 132552 65356
rect 131212 16584 131264 16590
rect 132512 16574 132540 65350
rect 132880 64530 132908 75958
rect 132972 69766 133000 79750
rect 133144 79688 133196 79694
rect 133144 79630 133196 79636
rect 133156 76498 133184 79630
rect 133328 79416 133380 79422
rect 133328 79358 133380 79364
rect 133340 78810 133368 79358
rect 133328 78804 133380 78810
rect 133328 78746 133380 78752
rect 133144 76492 133196 76498
rect 133144 76434 133196 76440
rect 133432 70394 133460 79784
rect 133558 79766 133610 79772
rect 133650 79824 133702 79830
rect 133650 79766 133702 79772
rect 133754 79778 133782 80036
rect 133846 79898 133874 80036
rect 133938 79966 133966 80036
rect 133926 79960 133978 79966
rect 134030 79937 134058 80036
rect 134122 79966 134150 80036
rect 134110 79960 134162 79966
rect 133926 79902 133978 79908
rect 134016 79928 134072 79937
rect 133834 79892 133886 79898
rect 134110 79902 134162 79908
rect 134016 79863 134072 79872
rect 133834 79834 133886 79840
rect 134214 79830 134242 80036
rect 134306 79898 134334 80036
rect 134398 79937 134426 80036
rect 134490 79966 134518 80036
rect 134478 79960 134530 79966
rect 134384 79928 134440 79937
rect 134294 79892 134346 79898
rect 134478 79902 134530 79908
rect 134384 79863 134440 79872
rect 134294 79834 134346 79840
rect 133972 79824 134024 79830
rect 133754 79750 133828 79778
rect 134202 79824 134254 79830
rect 134024 79784 134104 79812
rect 133972 79766 134024 79772
rect 133512 79688 133564 79694
rect 133512 79630 133564 79636
rect 133696 79688 133748 79694
rect 133696 79630 133748 79636
rect 133524 74225 133552 79630
rect 133708 78198 133736 79630
rect 133800 79608 133828 79750
rect 133800 79580 133920 79608
rect 133788 79416 133840 79422
rect 133788 79358 133840 79364
rect 133696 78192 133748 78198
rect 133696 78134 133748 78140
rect 133510 74216 133566 74225
rect 133510 74151 133566 74160
rect 133708 71126 133736 78134
rect 133800 72418 133828 79358
rect 133892 76022 133920 79580
rect 134076 76022 134104 79784
rect 134202 79766 134254 79772
rect 134338 79792 134394 79801
rect 134582 79744 134610 80036
rect 134674 79971 134702 80036
rect 134660 79962 134716 79971
rect 134660 79897 134716 79906
rect 134662 79824 134714 79830
rect 134338 79727 134394 79736
rect 134156 79688 134208 79694
rect 134156 79630 134208 79636
rect 134168 77382 134196 79630
rect 134248 79484 134300 79490
rect 134248 79426 134300 79432
rect 134260 78062 134288 79426
rect 134248 78056 134300 78062
rect 134248 77998 134300 78004
rect 134156 77376 134208 77382
rect 134156 77318 134208 77324
rect 133880 76016 133932 76022
rect 133880 75958 133932 75964
rect 134064 76016 134116 76022
rect 134064 75958 134116 75964
rect 134248 75268 134300 75274
rect 134248 75210 134300 75216
rect 134156 75064 134208 75070
rect 134156 75006 134208 75012
rect 133788 72412 133840 72418
rect 133788 72354 133840 72360
rect 133696 71120 133748 71126
rect 133696 71062 133748 71068
rect 133064 70366 133460 70394
rect 132960 69760 133012 69766
rect 132960 69702 133012 69708
rect 133064 65822 133092 70366
rect 133052 65816 133104 65822
rect 133052 65758 133104 65764
rect 133064 64874 133092 65758
rect 134168 65686 134196 75006
rect 134156 65680 134208 65686
rect 134156 65622 134208 65628
rect 134168 65414 134196 65622
rect 134156 65408 134208 65414
rect 134156 65350 134208 65356
rect 133064 64846 133184 64874
rect 132868 64524 132920 64530
rect 132868 64466 132920 64472
rect 133156 29646 133184 64846
rect 133788 64524 133840 64530
rect 133788 64466 133840 64472
rect 133800 55894 133828 64466
rect 134260 63306 134288 75210
rect 134352 66842 134380 79727
rect 134536 79716 134610 79744
rect 134660 79792 134662 79801
rect 134714 79792 134716 79801
rect 134660 79727 134716 79736
rect 134432 79688 134484 79694
rect 134432 79630 134484 79636
rect 134444 79286 134472 79630
rect 134432 79280 134484 79286
rect 134432 79222 134484 79228
rect 134432 76016 134484 76022
rect 134432 75958 134484 75964
rect 134340 66836 134392 66842
rect 134340 66778 134392 66784
rect 134248 63300 134300 63306
rect 134248 63242 134300 63248
rect 134260 62150 134288 63242
rect 134248 62144 134300 62150
rect 134248 62086 134300 62092
rect 133788 55888 133840 55894
rect 133788 55830 133840 55836
rect 134352 55214 134380 66778
rect 134444 64874 134472 75958
rect 134536 75070 134564 79716
rect 134766 79676 134794 80036
rect 134858 79830 134886 80036
rect 134846 79824 134898 79830
rect 134950 79801 134978 80036
rect 135042 79830 135070 80036
rect 135134 79937 135162 80036
rect 135120 79928 135176 79937
rect 135120 79863 135176 79872
rect 135226 79830 135254 80036
rect 135030 79824 135082 79830
rect 134846 79766 134898 79772
rect 134936 79792 134992 79801
rect 135030 79766 135082 79772
rect 135214 79824 135266 79830
rect 135318 79801 135346 80036
rect 135410 79966 135438 80036
rect 135502 79966 135530 80036
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135490 79960 135542 79966
rect 135490 79902 135542 79908
rect 135594 79812 135622 80036
rect 135686 79966 135714 80036
rect 135674 79960 135726 79966
rect 135674 79902 135726 79908
rect 135778 79812 135806 80036
rect 135870 79937 135898 80036
rect 135962 79966 135990 80036
rect 135950 79960 136002 79966
rect 135856 79928 135912 79937
rect 135950 79902 136002 79908
rect 135856 79863 135912 79872
rect 135214 79766 135266 79772
rect 135304 79792 135360 79801
rect 134936 79727 134992 79736
rect 135304 79727 135360 79736
rect 135456 79784 135622 79812
rect 135732 79784 135806 79812
rect 135904 79824 135956 79830
rect 135902 79792 135904 79801
rect 136054 79812 136082 80036
rect 136146 79966 136174 80036
rect 136238 79966 136266 80036
rect 136330 79966 136358 80036
rect 136422 79971 136450 80036
rect 136134 79960 136186 79966
rect 136134 79902 136186 79908
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 136408 79962 136464 79971
rect 136514 79966 136542 80036
rect 136408 79897 136464 79906
rect 136502 79960 136554 79966
rect 136502 79902 136554 79908
rect 136606 79835 136634 80036
rect 136698 79971 136726 80036
rect 136684 79962 136740 79971
rect 136684 79897 136740 79906
rect 136592 79826 136648 79835
rect 135956 79792 135958 79801
rect 135260 79688 135312 79694
rect 134766 79648 134840 79676
rect 134708 79552 134760 79558
rect 134708 79494 134760 79500
rect 134614 78568 134670 78577
rect 134614 78503 134670 78512
rect 134628 78169 134656 78503
rect 134614 78160 134670 78169
rect 134614 78095 134670 78104
rect 134524 75064 134576 75070
rect 134524 75006 134576 75012
rect 134628 68338 134656 78095
rect 134720 71774 134748 79494
rect 134812 75274 134840 79648
rect 135260 79630 135312 79636
rect 135352 79688 135404 79694
rect 135352 79630 135404 79636
rect 134984 79620 135036 79626
rect 134984 79562 135036 79568
rect 134892 79484 134944 79490
rect 134892 79426 134944 79432
rect 134904 78033 134932 79426
rect 134890 78024 134946 78033
rect 134890 77959 134946 77968
rect 134892 77376 134944 77382
rect 134892 77318 134944 77324
rect 134800 75268 134852 75274
rect 134800 75210 134852 75216
rect 134720 71746 134840 71774
rect 134616 68332 134668 68338
rect 134616 68274 134668 68280
rect 134708 65408 134760 65414
rect 134708 65350 134760 65356
rect 134444 64846 134656 64874
rect 134628 64666 134656 64846
rect 134616 64660 134668 64666
rect 134616 64602 134668 64608
rect 134352 55186 134564 55214
rect 133144 29640 133196 29646
rect 133144 29582 133196 29588
rect 132512 16546 133368 16574
rect 131212 16526 131264 16532
rect 130384 12436 130436 12442
rect 130384 12378 130436 12384
rect 133340 480 133368 16546
rect 134536 8974 134564 55186
rect 134628 18630 134656 64602
rect 134720 42158 134748 65350
rect 134812 64569 134840 71746
rect 134904 65958 134932 77318
rect 134996 72486 135024 79562
rect 135074 78432 135130 78441
rect 135074 78367 135130 78376
rect 135088 77722 135116 78367
rect 135076 77716 135128 77722
rect 135076 77658 135128 77664
rect 135272 75546 135300 79630
rect 135364 76090 135392 79630
rect 135456 78266 135484 79784
rect 135628 79688 135680 79694
rect 135628 79630 135680 79636
rect 135640 79121 135668 79630
rect 135732 79234 135760 79784
rect 136054 79784 136128 79812
rect 135902 79727 135958 79736
rect 135996 79688 136048 79694
rect 135996 79630 136048 79636
rect 135904 79620 135956 79626
rect 135904 79562 135956 79568
rect 135732 79206 135852 79234
rect 135626 79112 135682 79121
rect 135626 79047 135682 79056
rect 135824 78674 135852 79206
rect 135812 78668 135864 78674
rect 135812 78610 135864 78616
rect 135444 78260 135496 78266
rect 135444 78202 135496 78208
rect 135916 78180 135944 79562
rect 135732 78152 135944 78180
rect 135732 77217 135760 78152
rect 136008 78112 136036 79630
rect 135824 78084 136036 78112
rect 135718 77208 135774 77217
rect 135718 77143 135774 77152
rect 135628 76628 135680 76634
rect 135628 76570 135680 76576
rect 135536 76560 135588 76566
rect 135536 76502 135588 76508
rect 135352 76084 135404 76090
rect 135352 76026 135404 76032
rect 135260 75540 135312 75546
rect 135260 75482 135312 75488
rect 134984 72480 135036 72486
rect 134984 72422 135036 72428
rect 135548 68066 135576 76502
rect 135640 68406 135668 76570
rect 135720 76220 135772 76226
rect 135720 76162 135772 76168
rect 135628 68400 135680 68406
rect 135628 68342 135680 68348
rect 135536 68060 135588 68066
rect 135536 68002 135588 68008
rect 135444 67380 135496 67386
rect 135444 67322 135496 67328
rect 135260 67312 135312 67318
rect 135260 67254 135312 67260
rect 135272 66978 135300 67254
rect 135168 66972 135220 66978
rect 135168 66914 135220 66920
rect 135260 66972 135312 66978
rect 135260 66914 135312 66920
rect 135180 66638 135208 66914
rect 135456 66706 135484 67322
rect 135444 66700 135496 66706
rect 135444 66642 135496 66648
rect 135168 66632 135220 66638
rect 135168 66574 135220 66580
rect 134892 65952 134944 65958
rect 134892 65894 134944 65900
rect 134904 65686 134932 65894
rect 134892 65680 134944 65686
rect 134892 65622 134944 65628
rect 134798 64560 134854 64569
rect 134798 64495 134854 64504
rect 134812 63889 134840 64495
rect 134798 63880 134854 63889
rect 134798 63815 134854 63824
rect 134800 62144 134852 62150
rect 134800 62086 134852 62092
rect 134812 46238 134840 62086
rect 134800 46232 134852 46238
rect 134800 46174 134852 46180
rect 134708 42152 134760 42158
rect 134708 42094 134760 42100
rect 134616 18624 134668 18630
rect 134616 18566 134668 18572
rect 134524 8968 134576 8974
rect 134524 8910 134576 8916
rect 135456 3466 135484 66642
rect 135732 55214 135760 76162
rect 135824 68921 135852 78084
rect 135904 77988 135956 77994
rect 135904 77930 135956 77936
rect 135916 70281 135944 77930
rect 136100 76634 136128 79784
rect 136790 79778 136818 80036
rect 136882 79966 136910 80036
rect 136974 79971 137002 80036
rect 136870 79960 136922 79966
rect 136870 79902 136922 79908
rect 136960 79962 137016 79971
rect 137066 79966 137094 80036
rect 136960 79897 137016 79906
rect 137054 79960 137106 79966
rect 137054 79902 137106 79908
rect 137158 79898 137186 80036
rect 137146 79892 137198 79898
rect 137146 79834 137198 79840
rect 136180 79756 136232 79762
rect 136592 79761 136648 79770
rect 136180 79698 136232 79704
rect 136744 79750 136818 79778
rect 137100 79756 137152 79762
rect 136088 76628 136140 76634
rect 136088 76570 136140 76576
rect 136192 76158 136220 79698
rect 136456 79688 136508 79694
rect 136744 79642 136772 79750
rect 137250 79744 137278 80036
rect 137342 79971 137370 80036
rect 137328 79962 137384 79971
rect 137328 79897 137384 79906
rect 137434 79744 137462 80036
rect 137526 79971 137554 80036
rect 137512 79962 137568 79971
rect 137618 79966 137646 80036
rect 137710 79971 137738 80036
rect 137512 79897 137568 79906
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137696 79962 137752 79971
rect 137802 79966 137830 80036
rect 137894 79966 137922 80036
rect 137696 79897 137752 79906
rect 137790 79960 137842 79966
rect 137790 79902 137842 79908
rect 137882 79960 137934 79966
rect 137882 79902 137934 79908
rect 137986 79903 138014 80036
rect 138078 79966 138106 80036
rect 138170 79966 138198 80036
rect 138262 79971 138290 80036
rect 138066 79960 138118 79966
rect 137972 79894 138028 79903
rect 138066 79902 138118 79908
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 138248 79962 138304 79971
rect 138248 79897 138304 79906
rect 138354 79898 138382 80036
rect 138446 79971 138474 80036
rect 138432 79962 138488 79971
rect 137972 79829 138028 79838
rect 138342 79892 138394 79898
rect 138432 79897 138488 79906
rect 138538 79898 138566 80036
rect 138630 79971 138658 80036
rect 138616 79962 138672 79971
rect 138722 79966 138750 80036
rect 138342 79834 138394 79840
rect 138526 79892 138578 79898
rect 138616 79897 138672 79906
rect 138710 79960 138762 79966
rect 138710 79902 138762 79908
rect 138814 79898 138842 80036
rect 138906 79898 138934 80036
rect 138998 79966 139026 80036
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 138526 79834 138578 79840
rect 138802 79892 138854 79898
rect 138802 79834 138854 79840
rect 138894 79892 138946 79898
rect 138894 79834 138946 79840
rect 139090 79830 139118 80036
rect 138112 79824 138164 79830
rect 137250 79716 137324 79744
rect 137100 79698 137152 79704
rect 136456 79630 136508 79636
rect 136364 79620 136416 79626
rect 136364 79562 136416 79568
rect 136376 76566 136404 79562
rect 136364 76560 136416 76566
rect 136364 76502 136416 76508
rect 136468 76226 136496 79630
rect 136652 79614 136772 79642
rect 136916 79620 136968 79626
rect 136652 79121 136680 79614
rect 136916 79562 136968 79568
rect 137008 79620 137060 79626
rect 137008 79562 137060 79568
rect 136732 79552 136784 79558
rect 136732 79494 136784 79500
rect 136638 79112 136694 79121
rect 136638 79047 136694 79056
rect 136640 78668 136692 78674
rect 136640 78610 136692 78616
rect 136652 76809 136680 78610
rect 136744 78470 136772 79494
rect 136732 78464 136784 78470
rect 136732 78406 136784 78412
rect 136732 78056 136784 78062
rect 136732 77998 136784 78004
rect 136638 76800 136694 76809
rect 136638 76735 136694 76744
rect 136456 76220 136508 76226
rect 136456 76162 136508 76168
rect 136180 76152 136232 76158
rect 136086 76120 136142 76129
rect 136180 76094 136232 76100
rect 136548 76152 136600 76158
rect 136548 76094 136600 76100
rect 136086 76055 136142 76064
rect 136456 76084 136508 76090
rect 135902 70272 135958 70281
rect 135902 70207 135958 70216
rect 135810 68912 135866 68921
rect 135810 68847 135866 68856
rect 136100 67386 136128 76055
rect 136456 76026 136508 76032
rect 136362 75984 136418 75993
rect 136362 75919 136418 75928
rect 136376 68610 136404 75919
rect 136364 68604 136416 68610
rect 136364 68546 136416 68552
rect 136088 67380 136140 67386
rect 136088 67322 136140 67328
rect 136468 65890 136496 76026
rect 136560 70922 136588 76094
rect 136744 75177 136772 77998
rect 136824 76084 136876 76090
rect 136824 76026 136876 76032
rect 136730 75168 136786 75177
rect 136730 75103 136786 75112
rect 136548 70916 136600 70922
rect 136548 70858 136600 70864
rect 136456 65884 136508 65890
rect 136456 65826 136508 65832
rect 135904 65680 135956 65686
rect 135904 65622 135956 65628
rect 135720 55208 135772 55214
rect 135720 55150 135772 55156
rect 135916 3534 135944 65622
rect 136836 64462 136864 76026
rect 136928 66201 136956 79562
rect 137020 78810 137048 79562
rect 137008 78804 137060 78810
rect 137008 78746 137060 78752
rect 137020 77602 137048 78746
rect 137112 77761 137140 79698
rect 137190 79656 137246 79665
rect 137190 79591 137246 79600
rect 137098 77752 137154 77761
rect 137098 77687 137154 77696
rect 137020 77574 137140 77602
rect 137008 75268 137060 75274
rect 137008 75210 137060 75216
rect 137020 67386 137048 75210
rect 137008 67380 137060 67386
rect 137008 67322 137060 67328
rect 136914 66192 136970 66201
rect 136914 66127 136970 66136
rect 136824 64456 136876 64462
rect 136824 64398 136876 64404
rect 136836 64190 136864 64398
rect 136824 64184 136876 64190
rect 136824 64126 136876 64132
rect 137112 37942 137140 77574
rect 137204 67114 137232 79591
rect 137296 76090 137324 79716
rect 137388 79716 137462 79744
rect 137650 79792 137706 79801
rect 139078 79824 139130 79830
rect 138112 79766 138164 79772
rect 138294 79792 138350 79801
rect 137650 79727 137706 79736
rect 137388 79257 137416 79716
rect 137468 79620 137520 79626
rect 137468 79562 137520 79568
rect 137374 79248 137430 79257
rect 137374 79183 137430 79192
rect 137480 78985 137508 79562
rect 137466 78976 137522 78985
rect 137466 78911 137522 78920
rect 137376 77920 137428 77926
rect 137376 77862 137428 77868
rect 137284 76084 137336 76090
rect 137284 76026 137336 76032
rect 137388 69630 137416 77862
rect 137664 75274 137692 79727
rect 137742 79656 137798 79665
rect 137742 79591 137798 79600
rect 137836 79620 137888 79626
rect 137756 77625 137784 79591
rect 137836 79562 137888 79568
rect 137928 79620 137980 79626
rect 137928 79562 137980 79568
rect 138020 79620 138072 79626
rect 138020 79562 138072 79568
rect 137742 77616 137798 77625
rect 137742 77551 137798 77560
rect 137652 75268 137704 75274
rect 137652 75210 137704 75216
rect 137848 70394 137876 79562
rect 137940 77858 137968 79562
rect 138032 78742 138060 79562
rect 138020 78736 138072 78742
rect 138020 78678 138072 78684
rect 137928 77852 137980 77858
rect 137928 77794 137980 77800
rect 138020 76084 138072 76090
rect 138020 76026 138072 76032
rect 137848 70366 137968 70394
rect 137376 69624 137428 69630
rect 137376 69566 137428 69572
rect 137284 67380 137336 67386
rect 137284 67322 137336 67328
rect 137192 67108 137244 67114
rect 137192 67050 137244 67056
rect 137296 67046 137324 67322
rect 137284 67040 137336 67046
rect 137284 66982 137336 66988
rect 137296 47598 137324 66982
rect 137940 64874 137968 70366
rect 138032 67318 138060 76026
rect 138124 71774 138152 79766
rect 139182 79801 139210 80036
rect 139274 79937 139302 80036
rect 139260 79928 139316 79937
rect 139260 79863 139316 79872
rect 139366 79812 139394 80036
rect 139458 79937 139486 80036
rect 139550 79966 139578 80036
rect 139538 79960 139590 79966
rect 139444 79928 139500 79937
rect 139538 79902 139590 79908
rect 139444 79863 139500 79872
rect 139320 79801 139394 79812
rect 139078 79766 139130 79772
rect 139168 79792 139224 79801
rect 138294 79727 138350 79736
rect 138756 79756 138808 79762
rect 138124 71746 138244 71774
rect 138020 67312 138072 67318
rect 138020 67254 138072 67260
rect 138032 67114 138060 67254
rect 138020 67108 138072 67114
rect 138020 67050 138072 67056
rect 138216 65754 138244 71746
rect 138308 70394 138336 79727
rect 138756 79698 138808 79704
rect 138940 79756 138992 79762
rect 139168 79727 139224 79736
rect 139306 79792 139394 79801
rect 139362 79784 139394 79792
rect 139642 79778 139670 80036
rect 139734 79971 139762 80036
rect 139720 79962 139776 79971
rect 139720 79897 139776 79906
rect 139306 79727 139362 79736
rect 139492 79756 139544 79762
rect 138940 79698 138992 79704
rect 139492 79698 139544 79704
rect 139596 79750 139670 79778
rect 138572 79688 138624 79694
rect 138478 79656 138534 79665
rect 138572 79630 138624 79636
rect 138662 79656 138718 79665
rect 138478 79591 138534 79600
rect 138386 79384 138442 79393
rect 138386 79319 138442 79328
rect 138400 78606 138428 79319
rect 138388 78600 138440 78606
rect 138388 78542 138440 78548
rect 138388 77852 138440 77858
rect 138388 77794 138440 77800
rect 138400 71774 138428 77794
rect 138492 76022 138520 79591
rect 138584 77858 138612 79630
rect 138662 79591 138718 79600
rect 138572 77852 138624 77858
rect 138572 77794 138624 77800
rect 138572 77648 138624 77654
rect 138572 77590 138624 77596
rect 138480 76016 138532 76022
rect 138480 75958 138532 75964
rect 138584 74746 138612 77590
rect 138676 76945 138704 79591
rect 138768 77625 138796 79698
rect 138848 79620 138900 79626
rect 138848 79562 138900 79568
rect 138860 77790 138888 79562
rect 138952 78402 138980 79698
rect 139032 79688 139084 79694
rect 139032 79630 139084 79636
rect 139400 79688 139452 79694
rect 139400 79630 139452 79636
rect 138940 78396 138992 78402
rect 138940 78338 138992 78344
rect 138940 78260 138992 78266
rect 138940 78202 138992 78208
rect 138848 77784 138900 77790
rect 138848 77726 138900 77732
rect 138754 77616 138810 77625
rect 138754 77551 138810 77560
rect 138756 77512 138808 77518
rect 138756 77454 138808 77460
rect 138662 76936 138718 76945
rect 138662 76871 138718 76880
rect 138584 74718 138704 74746
rect 138400 71746 138612 71774
rect 138308 70366 138428 70394
rect 138400 68134 138428 70366
rect 138388 68128 138440 68134
rect 138388 68070 138440 68076
rect 138204 65748 138256 65754
rect 138204 65690 138256 65696
rect 137848 64846 137968 64874
rect 137848 64258 137876 64846
rect 137836 64252 137888 64258
rect 137836 64194 137888 64200
rect 137848 61470 137876 64194
rect 137836 61464 137888 61470
rect 137836 61406 137888 61412
rect 138584 53786 138612 71746
rect 138676 68746 138704 74718
rect 138768 73030 138796 77454
rect 138952 77194 138980 78202
rect 138860 77166 138980 77194
rect 138756 73024 138808 73030
rect 138756 72966 138808 72972
rect 138664 68740 138716 68746
rect 138664 68682 138716 68688
rect 138860 67561 138888 77166
rect 139044 76090 139072 79630
rect 139122 79384 139178 79393
rect 139122 79319 139178 79328
rect 139136 77314 139164 79319
rect 139306 79248 139362 79257
rect 139306 79183 139362 79192
rect 139124 77308 139176 77314
rect 139124 77250 139176 77256
rect 139032 76084 139084 76090
rect 139032 76026 139084 76032
rect 139124 76016 139176 76022
rect 139124 75958 139176 75964
rect 138940 73092 138992 73098
rect 138940 73034 138992 73040
rect 138846 67552 138902 67561
rect 138846 67487 138902 67496
rect 138664 67380 138716 67386
rect 138664 67322 138716 67328
rect 138676 66978 138704 67322
rect 138756 67108 138808 67114
rect 138756 67050 138808 67056
rect 138664 66972 138716 66978
rect 138664 66914 138716 66920
rect 138572 53780 138624 53786
rect 138572 53722 138624 53728
rect 137284 47592 137336 47598
rect 137284 47534 137336 47540
rect 137100 37936 137152 37942
rect 137100 37878 137152 37884
rect 137192 10396 137244 10402
rect 137192 10338 137244 10344
rect 135904 3528 135956 3534
rect 135904 3470 135956 3476
rect 135444 3460 135496 3466
rect 135444 3402 135496 3408
rect 137204 480 137232 10338
rect 138676 3466 138704 66914
rect 138768 22778 138796 67050
rect 138848 62144 138900 62150
rect 138848 62086 138900 62092
rect 138756 22772 138808 22778
rect 138756 22714 138808 22720
rect 138860 21418 138888 62086
rect 138952 52426 138980 73034
rect 139136 63442 139164 75958
rect 139320 67386 139348 79183
rect 139412 74497 139440 79630
rect 139504 79370 139532 79698
rect 139596 79472 139624 79750
rect 139826 79744 139854 80036
rect 139918 79966 139946 80036
rect 140010 79966 140038 80036
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139998 79960 140050 79966
rect 140102 79937 140130 80036
rect 139998 79902 140050 79908
rect 140088 79928 140144 79937
rect 140088 79863 140144 79872
rect 140044 79824 140096 79830
rect 139780 79716 139854 79744
rect 139950 79792 140006 79801
rect 140194 79812 140222 80036
rect 140286 79971 140314 80036
rect 140272 79962 140328 79971
rect 140272 79897 140328 79906
rect 140044 79766 140096 79772
rect 140148 79784 140222 79812
rect 139950 79727 140006 79736
rect 139596 79444 139716 79472
rect 139504 79342 139624 79370
rect 139492 79280 139544 79286
rect 139492 79222 139544 79228
rect 139398 74488 139454 74497
rect 139398 74423 139454 74432
rect 139504 68678 139532 79222
rect 139596 78878 139624 79342
rect 139584 78872 139636 78878
rect 139584 78814 139636 78820
rect 139688 78674 139716 79444
rect 139596 78646 139716 78674
rect 139596 76634 139624 78646
rect 139584 76628 139636 76634
rect 139584 76570 139636 76576
rect 139582 76392 139638 76401
rect 139582 76327 139638 76336
rect 139492 68672 139544 68678
rect 139492 68614 139544 68620
rect 139308 67380 139360 67386
rect 139308 67322 139360 67328
rect 139400 67380 139452 67386
rect 139400 67322 139452 67328
rect 139412 66774 139440 67322
rect 139400 66768 139452 66774
rect 139400 66710 139452 66716
rect 139124 63436 139176 63442
rect 139124 63378 139176 63384
rect 139136 62150 139164 63378
rect 139124 62144 139176 62150
rect 139124 62086 139176 62092
rect 138940 52420 138992 52426
rect 138940 52362 138992 52368
rect 138848 21412 138900 21418
rect 138848 21354 138900 21360
rect 139412 20670 139440 66710
rect 139400 20664 139452 20670
rect 139400 20606 139452 20612
rect 138664 3460 138716 3466
rect 138664 3402 138716 3408
rect 139504 3398 139532 68614
rect 139596 65482 139624 76327
rect 139780 67017 139808 79716
rect 139964 77586 139992 79727
rect 140056 77897 140084 79766
rect 140148 79393 140176 79784
rect 140378 79744 140406 80036
rect 140470 79778 140498 80036
rect 140562 79898 140590 80036
rect 140654 79937 140682 80036
rect 140640 79928 140696 79937
rect 140550 79892 140602 79898
rect 140640 79863 140696 79872
rect 140550 79834 140602 79840
rect 140746 79778 140774 80036
rect 140838 79898 140866 80036
rect 140930 79937 140958 80036
rect 140916 79928 140972 79937
rect 140826 79892 140878 79898
rect 140916 79863 140972 79872
rect 140826 79834 140878 79840
rect 141022 79812 141050 80036
rect 141114 79966 141142 80036
rect 141102 79960 141154 79966
rect 141102 79902 141154 79908
rect 141206 79898 141234 80036
rect 141298 79898 141326 80036
rect 141194 79892 141246 79898
rect 141194 79834 141246 79840
rect 141286 79892 141338 79898
rect 141286 79834 141338 79840
rect 140470 79750 140590 79778
rect 140240 79716 140406 79744
rect 140134 79384 140190 79393
rect 140134 79319 140190 79328
rect 140042 77888 140098 77897
rect 140042 77823 140098 77832
rect 139952 77580 140004 77586
rect 139952 77522 140004 77528
rect 140240 77178 140268 79716
rect 140562 79642 140590 79750
rect 140412 79620 140464 79626
rect 140412 79562 140464 79568
rect 140516 79614 140590 79642
rect 140700 79750 140774 79778
rect 140976 79784 141050 79812
rect 140424 78520 140452 79562
rect 140516 79286 140544 79614
rect 140700 79472 140728 79750
rect 140780 79688 140832 79694
rect 140832 79648 140912 79676
rect 140780 79630 140832 79636
rect 140608 79444 140728 79472
rect 140778 79520 140834 79529
rect 140778 79455 140780 79464
rect 140504 79280 140556 79286
rect 140504 79222 140556 79228
rect 140504 78804 140556 78810
rect 140504 78746 140556 78752
rect 140332 78492 140452 78520
rect 140332 77654 140360 78492
rect 140412 78396 140464 78402
rect 140412 78338 140464 78344
rect 140320 77648 140372 77654
rect 140320 77590 140372 77596
rect 140044 77172 140096 77178
rect 140044 77114 140096 77120
rect 140228 77172 140280 77178
rect 140228 77114 140280 77120
rect 139860 76628 139912 76634
rect 139860 76570 139912 76576
rect 139872 68542 139900 76570
rect 139952 75472 140004 75478
rect 139952 75414 140004 75420
rect 139964 75274 139992 75414
rect 139952 75268 140004 75274
rect 139952 75210 140004 75216
rect 140056 70394 140084 77114
rect 140424 77110 140452 78338
rect 140516 77926 140544 78746
rect 140504 77920 140556 77926
rect 140504 77862 140556 77868
rect 140608 77704 140636 79444
rect 140832 79455 140834 79464
rect 140780 79426 140832 79432
rect 140686 79384 140742 79393
rect 140686 79319 140742 79328
rect 140780 79348 140832 79354
rect 140516 77676 140636 77704
rect 140412 77104 140464 77110
rect 140412 77046 140464 77052
rect 140226 76800 140282 76809
rect 140226 76735 140282 76744
rect 139964 70366 140084 70394
rect 139860 68536 139912 68542
rect 139860 68478 139912 68484
rect 139766 67008 139822 67017
rect 139766 66943 139822 66952
rect 139584 65476 139636 65482
rect 139584 65418 139636 65424
rect 139964 60722 139992 70366
rect 140240 64954 140268 76735
rect 140516 67386 140544 77676
rect 140596 77580 140648 77586
rect 140596 77522 140648 77528
rect 140608 70990 140636 77522
rect 140596 70984 140648 70990
rect 140596 70926 140648 70932
rect 140504 67380 140556 67386
rect 140504 67322 140556 67328
rect 140700 66638 140728 79319
rect 140780 79290 140832 79296
rect 140792 79257 140820 79290
rect 140778 79248 140834 79257
rect 140778 79183 140834 79192
rect 140884 76106 140912 79648
rect 140976 76226 141004 79784
rect 141390 79778 141418 80036
rect 141482 79830 141510 80036
rect 141574 79830 141602 80036
rect 141666 79966 141694 80036
rect 141654 79960 141706 79966
rect 141654 79902 141706 79908
rect 141148 79756 141200 79762
rect 141148 79698 141200 79704
rect 141252 79750 141418 79778
rect 141470 79824 141522 79830
rect 141470 79766 141522 79772
rect 141562 79824 141614 79830
rect 141758 79778 141786 80036
rect 141850 79898 141878 80036
rect 141942 79966 141970 80036
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 141838 79892 141890 79898
rect 141838 79834 141890 79840
rect 142034 79778 142062 80036
rect 142126 79966 142154 80036
rect 142114 79960 142166 79966
rect 142114 79902 142166 79908
rect 142218 79812 142246 80036
rect 141562 79766 141614 79772
rect 141712 79750 141786 79778
rect 141884 79756 141936 79762
rect 141056 79688 141108 79694
rect 141056 79630 141108 79636
rect 141068 76498 141096 79630
rect 141056 76492 141108 76498
rect 141056 76434 141108 76440
rect 140964 76220 141016 76226
rect 140964 76162 141016 76168
rect 140884 76078 141004 76106
rect 140872 75336 140924 75342
rect 140872 75278 140924 75284
rect 140688 66632 140740 66638
rect 140688 66574 140740 66580
rect 140056 64926 140268 64954
rect 140056 64598 140084 64926
rect 140700 64874 140728 66574
rect 140884 65793 140912 75278
rect 140976 66065 141004 76078
rect 141056 75132 141108 75138
rect 141056 75074 141108 75080
rect 141068 67590 141096 75074
rect 141056 67584 141108 67590
rect 141056 67526 141108 67532
rect 141160 66230 141188 79698
rect 141252 79529 141280 79750
rect 141332 79688 141384 79694
rect 141424 79688 141476 79694
rect 141332 79630 141384 79636
rect 141422 79656 141424 79665
rect 141516 79688 141568 79694
rect 141476 79656 141478 79665
rect 141238 79520 141294 79529
rect 141238 79455 141294 79464
rect 141240 79348 141292 79354
rect 141240 79290 141292 79296
rect 141252 79257 141280 79290
rect 141238 79248 141294 79257
rect 141238 79183 141294 79192
rect 141238 78160 141294 78169
rect 141238 78095 141294 78104
rect 141252 68950 141280 78095
rect 141344 76634 141372 79630
rect 141516 79630 141568 79636
rect 141608 79688 141660 79694
rect 141608 79630 141660 79636
rect 141422 79591 141478 79600
rect 141424 79416 141476 79422
rect 141424 79358 141476 79364
rect 141436 79286 141464 79358
rect 141424 79280 141476 79286
rect 141424 79222 141476 79228
rect 141528 78538 141556 79630
rect 141516 78532 141568 78538
rect 141516 78474 141568 78480
rect 141424 77852 141476 77858
rect 141424 77794 141476 77800
rect 141332 76628 141384 76634
rect 141332 76570 141384 76576
rect 141240 68944 141292 68950
rect 141240 68886 141292 68892
rect 141436 68474 141464 77794
rect 141620 76616 141648 79630
rect 141712 77110 141740 79750
rect 141884 79698 141936 79704
rect 141988 79750 142062 79778
rect 142172 79784 142246 79812
rect 141700 77104 141752 77110
rect 141700 77046 141752 77052
rect 141528 76588 141648 76616
rect 141700 76628 141752 76634
rect 141528 68649 141556 76588
rect 141700 76570 141752 76576
rect 141608 76220 141660 76226
rect 141608 76162 141660 76168
rect 141620 68785 141648 76162
rect 141712 70009 141740 76570
rect 141792 76492 141844 76498
rect 141792 76434 141844 76440
rect 141698 70000 141754 70009
rect 141698 69935 141754 69944
rect 141606 68776 141662 68785
rect 141606 68711 141662 68720
rect 141514 68640 141570 68649
rect 141514 68575 141570 68584
rect 141424 68468 141476 68474
rect 141424 68410 141476 68416
rect 141148 66224 141200 66230
rect 141148 66166 141200 66172
rect 140962 66056 141018 66065
rect 140962 65991 141018 66000
rect 140870 65784 140926 65793
rect 140870 65719 140926 65728
rect 141804 64874 141832 76434
rect 141896 75138 141924 79698
rect 141988 75342 142016 79750
rect 141976 75336 142028 75342
rect 141976 75278 142028 75284
rect 141884 75132 141936 75138
rect 141884 75074 141936 75080
rect 142172 73914 142200 79784
rect 142310 79744 142338 80036
rect 142402 79966 142430 80036
rect 142494 79966 142522 80036
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142586 79830 142614 80036
rect 142574 79824 142626 79830
rect 142574 79766 142626 79772
rect 142678 79778 142706 80036
rect 142770 79898 142798 80036
rect 142758 79892 142810 79898
rect 142758 79834 142810 79840
rect 142862 79812 142890 80036
rect 142954 79937 142982 80036
rect 142940 79928 142996 79937
rect 142940 79863 142996 79872
rect 142862 79784 142936 79812
rect 142678 79750 142752 79778
rect 142724 79744 142752 79750
rect 142310 79716 142384 79744
rect 142724 79716 142798 79744
rect 142252 79620 142304 79626
rect 142252 79562 142304 79568
rect 142264 78266 142292 79562
rect 142356 79121 142384 79716
rect 142436 79688 142488 79694
rect 142436 79630 142488 79636
rect 142528 79688 142580 79694
rect 142528 79630 142580 79636
rect 142620 79688 142672 79694
rect 142770 79642 142798 79716
rect 142620 79630 142672 79636
rect 142342 79112 142398 79121
rect 142342 79047 142398 79056
rect 142344 78872 142396 78878
rect 142344 78814 142396 78820
rect 142252 78260 142304 78266
rect 142252 78202 142304 78208
rect 142356 77246 142384 78814
rect 142344 77240 142396 77246
rect 142344 77182 142396 77188
rect 142252 75472 142304 75478
rect 142252 75414 142304 75420
rect 142264 75274 142292 75414
rect 142344 75336 142396 75342
rect 142344 75278 142396 75284
rect 142252 75268 142304 75274
rect 142252 75210 142304 75216
rect 142160 73908 142212 73914
rect 142160 73850 142212 73856
rect 142066 70408 142122 70417
rect 142066 70343 142122 70352
rect 142080 68377 142108 70343
rect 142066 68368 142122 68377
rect 142066 68303 142122 68312
rect 142356 67250 142384 75278
rect 142448 75002 142476 79630
rect 142540 75070 142568 79630
rect 142632 78606 142660 79630
rect 142724 79614 142798 79642
rect 142620 78600 142672 78606
rect 142620 78542 142672 78548
rect 142620 76968 142672 76974
rect 142620 76910 142672 76916
rect 142632 76634 142660 76910
rect 142620 76628 142672 76634
rect 142620 76570 142672 76576
rect 142620 75268 142672 75274
rect 142620 75210 142672 75216
rect 142528 75064 142580 75070
rect 142528 75006 142580 75012
rect 142436 74996 142488 75002
rect 142436 74938 142488 74944
rect 142344 67244 142396 67250
rect 142344 67186 142396 67192
rect 142632 66230 142660 75210
rect 142620 66224 142672 66230
rect 142620 66166 142672 66172
rect 142724 66162 142752 79614
rect 142804 79552 142856 79558
rect 142804 79494 142856 79500
rect 142816 79121 142844 79494
rect 142802 79112 142858 79121
rect 142802 79047 142858 79056
rect 142804 78600 142856 78606
rect 142804 78542 142856 78548
rect 142816 75274 142844 78542
rect 142908 75342 142936 79784
rect 143046 79778 143074 80036
rect 143138 79966 143166 80036
rect 143126 79960 143178 79966
rect 143126 79902 143178 79908
rect 143230 79812 143258 80036
rect 143000 79750 143074 79778
rect 143184 79784 143258 79812
rect 143000 78878 143028 79750
rect 143080 79688 143132 79694
rect 143080 79630 143132 79636
rect 142988 78872 143040 78878
rect 142988 78814 143040 78820
rect 143092 78441 143120 79630
rect 143078 78432 143134 78441
rect 143078 78367 143134 78376
rect 143080 77104 143132 77110
rect 143080 77046 143132 77052
rect 142896 75336 142948 75342
rect 142896 75278 142948 75284
rect 142988 75336 143040 75342
rect 142988 75278 143040 75284
rect 142804 75268 142856 75274
rect 142804 75210 142856 75216
rect 143000 75070 143028 75278
rect 142988 75064 143040 75070
rect 142988 75006 143040 75012
rect 142804 74996 142856 75002
rect 142804 74938 142856 74944
rect 142816 69766 142844 74938
rect 142988 73024 143040 73030
rect 142988 72966 143040 72972
rect 143000 72622 143028 72966
rect 142988 72616 143040 72622
rect 142988 72558 143040 72564
rect 142804 69760 142856 69766
rect 142804 69702 142856 69708
rect 142804 67244 142856 67250
rect 142804 67186 142856 67192
rect 142712 66156 142764 66162
rect 142712 66098 142764 66104
rect 140148 64846 140728 64874
rect 141436 64846 141832 64874
rect 140044 64592 140096 64598
rect 140044 64534 140096 64540
rect 139952 60716 140004 60722
rect 139952 60658 140004 60664
rect 140056 43450 140084 64534
rect 140148 49026 140176 64846
rect 141436 63374 141464 64846
rect 141424 63368 141476 63374
rect 141424 63310 141476 63316
rect 141436 53174 141464 63310
rect 141424 53168 141476 53174
rect 141424 53110 141476 53116
rect 140136 49020 140188 49026
rect 140136 48962 140188 48968
rect 140044 43444 140096 43450
rect 140044 43386 140096 43392
rect 142816 10334 142844 67186
rect 142896 66224 142948 66230
rect 142896 66166 142948 66172
rect 142908 65278 142936 66166
rect 142896 65272 142948 65278
rect 142896 65214 142948 65220
rect 142908 13122 142936 65214
rect 143000 62830 143028 72558
rect 143092 63510 143120 77046
rect 143184 73030 143212 79784
rect 143322 79744 143350 80036
rect 143414 79966 143442 80036
rect 143506 79971 143534 80036
rect 143402 79960 143454 79966
rect 143402 79902 143454 79908
rect 143492 79962 143548 79971
rect 143492 79897 143548 79906
rect 143492 79792 143548 79801
rect 143276 79716 143350 79744
rect 143460 79736 143492 79744
rect 143598 79778 143626 80036
rect 143690 79898 143718 80036
rect 143782 79898 143810 80036
rect 143678 79892 143730 79898
rect 143678 79834 143730 79840
rect 143770 79892 143822 79898
rect 143770 79834 143822 79840
rect 143722 79792 143778 79801
rect 143598 79750 143722 79778
rect 143460 79727 143548 79736
rect 143874 79744 143902 80036
rect 143966 79898 143994 80036
rect 144058 79898 144086 80036
rect 144150 79966 144178 80036
rect 144242 79966 144270 80036
rect 144334 79966 144362 80036
rect 144138 79960 144190 79966
rect 144138 79902 144190 79908
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 143954 79892 144006 79898
rect 143954 79834 144006 79840
rect 144046 79892 144098 79898
rect 144046 79834 144098 79840
rect 144426 79812 144454 80036
rect 144518 79898 144546 80036
rect 144610 79898 144638 80036
rect 144506 79892 144558 79898
rect 144506 79834 144558 79840
rect 144598 79892 144650 79898
rect 144598 79834 144650 79840
rect 144274 79792 144330 79801
rect 144184 79756 144236 79762
rect 143722 79727 143778 79736
rect 143460 79716 143534 79727
rect 143828 79716 143902 79744
rect 144012 79716 144184 79744
rect 143276 78674 143304 79716
rect 143356 79620 143408 79626
rect 143356 79562 143408 79568
rect 143264 78668 143316 78674
rect 143264 78610 143316 78616
rect 143172 73024 143224 73030
rect 143172 72966 143224 72972
rect 143368 71738 143396 79562
rect 143460 78577 143488 79716
rect 143632 79688 143684 79694
rect 143828 79676 143856 79716
rect 143632 79630 143684 79636
rect 143736 79648 143856 79676
rect 143540 79552 143592 79558
rect 143540 79494 143592 79500
rect 143446 78568 143502 78577
rect 143446 78503 143502 78512
rect 143552 74440 143580 79494
rect 143460 74412 143580 74440
rect 143460 73658 143488 74412
rect 143540 74316 143592 74322
rect 143540 74258 143592 74264
rect 143552 73846 143580 74258
rect 143540 73840 143592 73846
rect 143540 73782 143592 73788
rect 143460 73630 143580 73658
rect 143356 71732 143408 71738
rect 143356 71674 143408 71680
rect 143368 70394 143396 71674
rect 143552 71330 143580 73630
rect 143644 73098 143672 79630
rect 143632 73092 143684 73098
rect 143632 73034 143684 73040
rect 143736 71738 143764 79648
rect 143908 79620 143960 79626
rect 143908 79562 143960 79568
rect 143816 79552 143868 79558
rect 143816 79494 143868 79500
rect 143828 72593 143856 79494
rect 143920 75274 143948 79562
rect 143908 75268 143960 75274
rect 143908 75210 143960 75216
rect 143814 72584 143870 72593
rect 143814 72519 143870 72528
rect 143724 71732 143776 71738
rect 143724 71674 143776 71680
rect 143736 71398 143764 71674
rect 143724 71392 143776 71398
rect 143724 71334 143776 71340
rect 143540 71324 143592 71330
rect 143540 71266 143592 71272
rect 143368 70366 143488 70394
rect 143460 69698 143488 70366
rect 143448 69692 143500 69698
rect 143448 69634 143500 69640
rect 144012 67522 144040 79716
rect 144274 79727 144330 79736
rect 144380 79784 144454 79812
rect 144184 79698 144236 79704
rect 144184 79620 144236 79626
rect 144184 79562 144236 79568
rect 144092 79552 144144 79558
rect 144092 79494 144144 79500
rect 144104 73098 144132 79494
rect 144196 73846 144224 79562
rect 144288 75426 144316 79727
rect 144380 78849 144408 79784
rect 144460 79688 144512 79694
rect 144460 79630 144512 79636
rect 144366 78840 144422 78849
rect 144366 78775 144422 78784
rect 144366 78160 144422 78169
rect 144366 78095 144422 78104
rect 144380 77858 144408 78095
rect 144472 77897 144500 79630
rect 144552 79620 144604 79626
rect 144702 79608 144730 80036
rect 144794 79937 144822 80036
rect 144886 79966 144914 80036
rect 144978 79966 145006 80036
rect 145070 79966 145098 80036
rect 145162 79966 145190 80036
rect 145254 79971 145282 80036
rect 144874 79960 144926 79966
rect 144780 79928 144836 79937
rect 144874 79902 144926 79908
rect 144966 79960 145018 79966
rect 144966 79902 145018 79908
rect 145058 79960 145110 79966
rect 145058 79902 145110 79908
rect 145150 79960 145202 79966
rect 145150 79902 145202 79908
rect 145240 79962 145296 79971
rect 145240 79897 145296 79906
rect 144780 79863 144836 79872
rect 144828 79824 144880 79830
rect 144828 79766 144880 79772
rect 145104 79824 145156 79830
rect 145104 79766 145156 79772
rect 145196 79824 145248 79830
rect 145346 79812 145374 80036
rect 145438 79966 145466 80036
rect 145426 79960 145478 79966
rect 145426 79902 145478 79908
rect 145346 79784 145420 79812
rect 145196 79766 145248 79772
rect 144840 79665 144868 79766
rect 144920 79756 144972 79762
rect 144920 79698 144972 79704
rect 144552 79562 144604 79568
rect 144656 79580 144730 79608
rect 144826 79656 144882 79665
rect 144826 79591 144882 79600
rect 144458 77888 144514 77897
rect 144368 77852 144420 77858
rect 144458 77823 144514 77832
rect 144368 77794 144420 77800
rect 144564 76537 144592 79562
rect 144656 78810 144684 79580
rect 144826 79520 144882 79529
rect 144826 79455 144882 79464
rect 144644 78804 144696 78810
rect 144644 78746 144696 78752
rect 144840 77586 144868 79455
rect 144932 79150 144960 79698
rect 145012 79688 145064 79694
rect 145116 79665 145144 79766
rect 145012 79630 145064 79636
rect 145102 79656 145158 79665
rect 144920 79144 144972 79150
rect 144920 79086 144972 79092
rect 145024 78554 145052 79630
rect 145102 79591 145158 79600
rect 145024 78526 145144 78554
rect 145010 78432 145066 78441
rect 145010 78367 145066 78376
rect 144828 77580 144880 77586
rect 144828 77522 144880 77528
rect 145024 76634 145052 78367
rect 145012 76628 145064 76634
rect 145012 76570 145064 76576
rect 144550 76528 144606 76537
rect 144550 76463 144606 76472
rect 144288 75398 144408 75426
rect 145116 75410 145144 78526
rect 144276 75268 144328 75274
rect 144276 75210 144328 75216
rect 144184 73840 144236 73846
rect 144184 73782 144236 73788
rect 144092 73092 144144 73098
rect 144092 73034 144144 73040
rect 144184 71732 144236 71738
rect 144184 71674 144236 71680
rect 144000 67516 144052 67522
rect 144000 67458 144052 67464
rect 143448 66156 143500 66162
rect 143448 66098 143500 66104
rect 143460 65550 143488 66098
rect 143448 65544 143500 65550
rect 143448 65486 143500 65492
rect 144012 64258 144040 67458
rect 144000 64252 144052 64258
rect 144000 64194 144052 64200
rect 143080 63504 143132 63510
rect 143080 63446 143132 63452
rect 142988 62824 143040 62830
rect 142988 62766 143040 62772
rect 144196 21486 144224 71674
rect 144288 67454 144316 75210
rect 144380 71262 144408 75398
rect 145104 75404 145156 75410
rect 145104 75346 145156 75352
rect 145208 75041 145236 79766
rect 145286 79656 145342 79665
rect 145286 79591 145342 79600
rect 145300 79286 145328 79591
rect 145288 79280 145340 79286
rect 145288 79222 145340 79228
rect 145288 79144 145340 79150
rect 145288 79086 145340 79092
rect 145194 75032 145250 75041
rect 145194 74967 145250 74976
rect 145300 73982 145328 79086
rect 145288 73976 145340 73982
rect 145288 73918 145340 73924
rect 145300 73154 145328 73918
rect 145208 73126 145328 73154
rect 144460 73092 144512 73098
rect 144460 73034 144512 73040
rect 144472 72690 144500 73034
rect 144460 72684 144512 72690
rect 144460 72626 144512 72632
rect 144368 71256 144420 71262
rect 144368 71198 144420 71204
rect 144276 67448 144328 67454
rect 144276 67390 144328 67396
rect 144288 28286 144316 67390
rect 144380 43518 144408 71198
rect 144472 60042 144500 72626
rect 145208 72486 145236 73126
rect 145196 72480 145248 72486
rect 145196 72422 145248 72428
rect 145392 70378 145420 79784
rect 145530 79744 145558 80036
rect 145622 79971 145650 80036
rect 145608 79962 145664 79971
rect 145608 79897 145664 79906
rect 145714 79898 145742 80036
rect 145806 79966 145834 80036
rect 145898 79971 145926 80036
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145884 79962 145940 79971
rect 145990 79966 146018 80036
rect 146082 79966 146110 80036
rect 146174 79971 146202 80036
rect 145702 79892 145754 79898
rect 145884 79897 145940 79906
rect 145978 79960 146030 79966
rect 145978 79902 146030 79908
rect 146070 79960 146122 79966
rect 146070 79902 146122 79908
rect 146160 79962 146216 79971
rect 146160 79897 146216 79906
rect 146266 79898 146294 80036
rect 146358 79903 146386 80036
rect 146450 79966 146478 80036
rect 146438 79960 146490 79966
rect 145702 79834 145754 79840
rect 146254 79892 146306 79898
rect 146254 79834 146306 79840
rect 146344 79894 146400 79903
rect 146438 79902 146490 79908
rect 146344 79829 146400 79838
rect 145484 79716 145558 79744
rect 145656 79756 145708 79762
rect 145484 79558 145512 79716
rect 145656 79698 145708 79704
rect 145748 79756 145800 79762
rect 145748 79698 145800 79704
rect 145932 79756 145984 79762
rect 145932 79698 145984 79704
rect 146116 79756 146168 79762
rect 146116 79698 146168 79704
rect 146208 79756 146260 79762
rect 146208 79698 146260 79704
rect 146392 79756 146444 79762
rect 146542 79744 146570 80036
rect 146634 79966 146662 80036
rect 146622 79960 146674 79966
rect 146622 79902 146674 79908
rect 146392 79698 146444 79704
rect 146496 79716 146570 79744
rect 145562 79656 145618 79665
rect 145562 79591 145564 79600
rect 145616 79591 145618 79600
rect 145564 79562 145616 79568
rect 145472 79552 145524 79558
rect 145472 79494 145524 79500
rect 145470 79384 145526 79393
rect 145470 79319 145526 79328
rect 145380 70372 145432 70378
rect 145380 70314 145432 70320
rect 145484 69902 145512 79319
rect 145564 79280 145616 79286
rect 145564 79222 145616 79228
rect 145576 72457 145604 79222
rect 145668 75857 145696 79698
rect 145760 79150 145788 79698
rect 145840 79552 145892 79558
rect 145840 79494 145892 79500
rect 145748 79144 145800 79150
rect 145748 79086 145800 79092
rect 145852 75914 145880 79494
rect 145760 75886 145880 75914
rect 145654 75848 145710 75857
rect 145654 75783 145710 75792
rect 145760 74118 145788 75886
rect 145944 75614 145972 79698
rect 146024 79688 146076 79694
rect 146024 79630 146076 79636
rect 146036 78033 146064 79630
rect 146128 79014 146156 79698
rect 146116 79008 146168 79014
rect 146116 78950 146168 78956
rect 146116 78804 146168 78810
rect 146116 78746 146168 78752
rect 146022 78024 146078 78033
rect 146022 77959 146078 77968
rect 146128 76906 146156 78746
rect 146116 76900 146168 76906
rect 146116 76842 146168 76848
rect 145932 75608 145984 75614
rect 145932 75550 145984 75556
rect 146220 75478 146248 79698
rect 146298 79656 146354 79665
rect 146298 79591 146354 79600
rect 146312 77518 146340 79591
rect 146300 77512 146352 77518
rect 146300 77454 146352 77460
rect 146208 75472 146260 75478
rect 146208 75414 146260 75420
rect 146404 75410 146432 79698
rect 146392 75404 146444 75410
rect 146392 75346 146444 75352
rect 145748 74112 145800 74118
rect 145748 74054 145800 74060
rect 145562 72448 145618 72457
rect 145562 72383 145618 72392
rect 145760 70394 145788 74054
rect 145564 70372 145616 70378
rect 145564 70314 145616 70320
rect 145668 70366 145788 70394
rect 145472 69896 145524 69902
rect 145472 69838 145524 69844
rect 144920 64184 144972 64190
rect 144920 64126 144972 64132
rect 144460 60036 144512 60042
rect 144460 59978 144512 59984
rect 144368 43512 144420 43518
rect 144368 43454 144420 43460
rect 144276 28280 144328 28286
rect 144276 28222 144328 28228
rect 144184 21480 144236 21486
rect 144184 21422 144236 21428
rect 142896 13116 142948 13122
rect 142896 13058 142948 13064
rect 142804 10328 142856 10334
rect 142804 10270 142856 10276
rect 141056 3528 141108 3534
rect 141056 3470 141108 3476
rect 139492 3392 139544 3398
rect 139492 3334 139544 3340
rect 141068 480 141096 3470
rect 144932 480 144960 64126
rect 145576 9042 145604 70314
rect 145668 54602 145696 70366
rect 146496 68202 146524 79716
rect 146726 79676 146754 80036
rect 146818 79898 146846 80036
rect 146910 79966 146938 80036
rect 146898 79960 146950 79966
rect 146898 79902 146950 79908
rect 146806 79892 146858 79898
rect 146806 79834 146858 79840
rect 147002 79812 147030 80036
rect 147094 79937 147122 80036
rect 147080 79928 147136 79937
rect 147080 79863 147136 79872
rect 147002 79784 147076 79812
rect 147048 79778 147076 79784
rect 147048 79750 147122 79778
rect 146588 79648 146754 79676
rect 146944 79688 146996 79694
rect 146588 68814 146616 79648
rect 146944 79630 146996 79636
rect 146668 79552 146720 79558
rect 146668 79494 146720 79500
rect 146758 79520 146814 79529
rect 146680 75546 146708 79494
rect 146758 79455 146814 79464
rect 146668 75540 146720 75546
rect 146668 75482 146720 75488
rect 146772 70394 146800 79455
rect 146852 75404 146904 75410
rect 146852 75346 146904 75352
rect 146680 70366 146800 70394
rect 146576 68808 146628 68814
rect 146576 68750 146628 68756
rect 146484 68196 146536 68202
rect 146484 68138 146536 68144
rect 146680 64802 146708 70366
rect 146864 70242 146892 75346
rect 146956 73817 146984 79630
rect 147094 79540 147122 79750
rect 147186 79744 147214 80036
rect 147278 79966 147306 80036
rect 147370 79966 147398 80036
rect 147462 79971 147490 80036
rect 147266 79960 147318 79966
rect 147266 79902 147318 79908
rect 147358 79960 147410 79966
rect 147358 79902 147410 79908
rect 147448 79962 147504 79971
rect 147554 79966 147582 80036
rect 147646 79971 147674 80036
rect 147448 79897 147504 79906
rect 147542 79960 147594 79966
rect 147542 79902 147594 79908
rect 147632 79962 147688 79971
rect 147738 79966 147766 80036
rect 147632 79897 147688 79906
rect 147726 79960 147778 79966
rect 147726 79902 147778 79908
rect 147312 79824 147364 79830
rect 147680 79824 147732 79830
rect 147312 79766 147364 79772
rect 147586 79792 147642 79801
rect 147186 79716 147260 79744
rect 147048 79512 147122 79540
rect 146942 73808 146998 73817
rect 146942 73743 146998 73752
rect 147048 71505 147076 79512
rect 147232 73154 147260 79716
rect 147324 78033 147352 79766
rect 147404 79756 147456 79762
rect 147830 79812 147858 80036
rect 147922 79898 147950 80036
rect 147910 79892 147962 79898
rect 147910 79834 147962 79840
rect 147680 79766 147732 79772
rect 147784 79784 147858 79812
rect 147586 79727 147642 79736
rect 147404 79698 147456 79704
rect 147416 78402 147444 79698
rect 147496 79688 147548 79694
rect 147496 79630 147548 79636
rect 147404 78396 147456 78402
rect 147404 78338 147456 78344
rect 147310 78024 147366 78033
rect 147310 77959 147366 77968
rect 147140 73126 147260 73154
rect 147034 71496 147090 71505
rect 147034 71431 147090 71440
rect 147036 71324 147088 71330
rect 147036 71266 147088 71272
rect 146852 70236 146904 70242
rect 146852 70178 146904 70184
rect 146944 65884 146996 65890
rect 146944 65826 146996 65832
rect 146668 64796 146720 64802
rect 146668 64738 146720 64744
rect 145656 54596 145708 54602
rect 145656 54538 145708 54544
rect 145564 9036 145616 9042
rect 145564 8978 145616 8984
rect 146956 3534 146984 65826
rect 147048 45558 147076 71266
rect 147140 67182 147168 73126
rect 147508 72350 147536 79630
rect 147600 76838 147628 79727
rect 147588 76832 147640 76838
rect 147588 76774 147640 76780
rect 147692 74254 147720 79766
rect 147784 77858 147812 79784
rect 148014 79778 148042 80036
rect 148106 79898 148134 80036
rect 148198 79898 148226 80036
rect 148094 79892 148146 79898
rect 148094 79834 148146 79840
rect 148186 79892 148238 79898
rect 148186 79834 148238 79840
rect 148290 79835 148318 80036
rect 147922 79750 148042 79778
rect 148276 79826 148332 79835
rect 148382 79830 148410 80036
rect 148474 79966 148502 80036
rect 148462 79960 148514 79966
rect 148566 79937 148594 80036
rect 148462 79902 148514 79908
rect 148552 79928 148608 79937
rect 148552 79863 148608 79872
rect 148276 79761 148332 79770
rect 148370 79824 148422 79830
rect 148658 79812 148686 80036
rect 148750 79966 148778 80036
rect 148738 79960 148790 79966
rect 148738 79902 148790 79908
rect 148842 79898 148870 80036
rect 148934 79966 148962 80036
rect 148922 79960 148974 79966
rect 148922 79902 148974 79908
rect 148830 79892 148882 79898
rect 148830 79834 148882 79840
rect 148658 79784 148778 79812
rect 148370 79766 148422 79772
rect 147922 79744 147950 79750
rect 148750 79744 148778 79784
rect 149026 79744 149054 80036
rect 149118 79937 149146 80036
rect 149210 79966 149238 80036
rect 149198 79960 149250 79966
rect 149104 79928 149160 79937
rect 149198 79902 149250 79908
rect 149104 79863 149160 79872
rect 147876 79716 147950 79744
rect 148704 79716 148778 79744
rect 148980 79716 149054 79744
rect 149302 79744 149330 80036
rect 149394 79966 149422 80036
rect 149486 79971 149514 80036
rect 149382 79960 149434 79966
rect 149382 79902 149434 79908
rect 149472 79962 149528 79971
rect 149472 79897 149528 79906
rect 149578 79898 149606 80036
rect 149670 79966 149698 80036
rect 149762 79971 149790 80036
rect 149658 79960 149710 79966
rect 149658 79902 149710 79908
rect 149748 79962 149804 79971
rect 149854 79966 149882 80036
rect 149946 79966 149974 80036
rect 149566 79892 149618 79898
rect 149748 79897 149804 79906
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149934 79960 149986 79966
rect 150038 79937 150066 80036
rect 149934 79902 149986 79908
rect 150024 79928 150080 79937
rect 150024 79863 150080 79872
rect 149566 79834 149618 79840
rect 149978 79792 150034 79801
rect 149302 79716 149376 79744
rect 149978 79727 150034 79736
rect 150130 79744 150158 80036
rect 150222 79903 150250 80036
rect 150208 79894 150264 79903
rect 150314 79898 150342 80036
rect 150406 79903 150434 80036
rect 150498 79966 150526 80036
rect 150486 79960 150538 79966
rect 150208 79829 150264 79838
rect 150302 79892 150354 79898
rect 150302 79834 150354 79840
rect 150392 79894 150448 79903
rect 150486 79902 150538 79908
rect 150392 79829 150448 79838
rect 150590 79812 150618 80036
rect 150682 79937 150710 80036
rect 150668 79928 150724 79937
rect 150774 79898 150802 80036
rect 150668 79863 150724 79872
rect 150762 79892 150814 79898
rect 150762 79834 150814 79840
rect 150544 79784 150618 79812
rect 150256 79756 150308 79762
rect 147772 77852 147824 77858
rect 147772 77794 147824 77800
rect 147772 77580 147824 77586
rect 147772 77522 147824 77528
rect 147784 74458 147812 77522
rect 147772 74452 147824 74458
rect 147772 74394 147824 74400
rect 147680 74248 147732 74254
rect 147680 74190 147732 74196
rect 147496 72344 147548 72350
rect 147496 72286 147548 72292
rect 147692 70394 147720 74190
rect 147876 72758 147904 79716
rect 148232 79688 148284 79694
rect 148046 79656 148102 79665
rect 147956 79620 148008 79626
rect 148046 79591 148102 79600
rect 148230 79656 148232 79665
rect 148508 79688 148560 79694
rect 148284 79656 148286 79665
rect 148508 79630 148560 79636
rect 148600 79688 148652 79694
rect 148600 79630 148652 79636
rect 148230 79591 148286 79600
rect 147956 79562 148008 79568
rect 147968 76673 147996 79562
rect 147954 76664 148010 76673
rect 147954 76599 148010 76608
rect 148060 73642 148088 79591
rect 148232 79552 148284 79558
rect 148232 79494 148284 79500
rect 148414 79520 148470 79529
rect 148140 75200 148192 75206
rect 148140 75142 148192 75148
rect 148048 73636 148100 73642
rect 148048 73578 148100 73584
rect 147864 72752 147916 72758
rect 147864 72694 147916 72700
rect 147692 70366 147812 70394
rect 147128 67176 147180 67182
rect 147128 67118 147180 67124
rect 147036 45552 147088 45558
rect 147036 45494 147088 45500
rect 147784 28966 147812 70366
rect 148152 66910 148180 75142
rect 148244 69834 148272 79494
rect 148414 79455 148470 79464
rect 148324 77988 148376 77994
rect 148324 77930 148376 77936
rect 148336 75206 148364 77930
rect 148428 75585 148456 79455
rect 148520 78810 148548 79630
rect 148508 78804 148560 78810
rect 148508 78746 148560 78752
rect 148612 78305 148640 79630
rect 148598 78296 148654 78305
rect 148598 78231 148654 78240
rect 148600 77852 148652 77858
rect 148600 77794 148652 77800
rect 148414 75576 148470 75585
rect 148414 75511 148470 75520
rect 148324 75200 148376 75206
rect 148324 75142 148376 75148
rect 148612 69970 148640 77794
rect 148704 77586 148732 79716
rect 148876 79688 148928 79694
rect 148796 79648 148876 79676
rect 148796 78130 148824 79648
rect 148980 79665 149008 79716
rect 148876 79630 148928 79636
rect 148966 79656 149022 79665
rect 149150 79656 149206 79665
rect 148966 79591 149022 79600
rect 149060 79620 149112 79626
rect 149150 79591 149206 79600
rect 149244 79620 149296 79626
rect 149060 79562 149112 79568
rect 148968 79552 149020 79558
rect 148968 79494 149020 79500
rect 148876 78260 148928 78266
rect 148876 78202 148928 78208
rect 148784 78124 148836 78130
rect 148784 78066 148836 78072
rect 148692 77580 148744 77586
rect 148692 77522 148744 77528
rect 148888 73710 148916 78202
rect 148980 77994 149008 79494
rect 149072 79014 149100 79562
rect 149060 79008 149112 79014
rect 149060 78950 149112 78956
rect 148968 77988 149020 77994
rect 148968 77930 149020 77936
rect 148876 73704 148928 73710
rect 148876 73646 148928 73652
rect 149164 71670 149192 79591
rect 149244 79562 149296 79568
rect 149256 76770 149284 79562
rect 149244 76764 149296 76770
rect 149244 76706 149296 76712
rect 149348 75914 149376 79716
rect 149428 79688 149480 79694
rect 149428 79630 149480 79636
rect 149612 79688 149664 79694
rect 149612 79630 149664 79636
rect 149440 78033 149468 79630
rect 149518 79384 149574 79393
rect 149518 79319 149574 79328
rect 149426 78024 149482 78033
rect 149426 77959 149482 77968
rect 149256 75886 149376 75914
rect 149256 75682 149284 75886
rect 149244 75676 149296 75682
rect 149244 75618 149296 75624
rect 149152 71664 149204 71670
rect 149152 71606 149204 71612
rect 149532 71194 149560 79319
rect 149624 76702 149652 79630
rect 149796 79620 149848 79626
rect 149796 79562 149848 79568
rect 149704 79552 149756 79558
rect 149704 79494 149756 79500
rect 149612 76696 149664 76702
rect 149612 76638 149664 76644
rect 149716 74934 149744 79494
rect 149704 74928 149756 74934
rect 149704 74870 149756 74876
rect 149808 71466 149836 79562
rect 149992 78334 150020 79727
rect 150130 79716 150204 79744
rect 149980 78328 150032 78334
rect 149980 78270 150032 78276
rect 150176 75886 150204 79716
rect 150256 79698 150308 79704
rect 150440 79756 150492 79762
rect 150440 79698 150492 79704
rect 150268 78033 150296 79698
rect 150346 79656 150402 79665
rect 150346 79591 150402 79600
rect 150360 79218 150388 79591
rect 150348 79212 150400 79218
rect 150348 79154 150400 79160
rect 150254 78024 150310 78033
rect 150254 77959 150310 77968
rect 150164 75880 150216 75886
rect 150164 75822 150216 75828
rect 150164 75676 150216 75682
rect 150164 75618 150216 75624
rect 149888 71664 149940 71670
rect 149888 71606 149940 71612
rect 149796 71460 149848 71466
rect 149796 71402 149848 71408
rect 149520 71188 149572 71194
rect 149520 71130 149572 71136
rect 149532 70394 149560 71130
rect 149532 70366 149744 70394
rect 148600 69964 148652 69970
rect 148600 69906 148652 69912
rect 148232 69828 148284 69834
rect 148232 69770 148284 69776
rect 148140 66904 148192 66910
rect 148140 66846 148192 66852
rect 148324 66904 148376 66910
rect 148324 66846 148376 66852
rect 148336 40730 148364 66846
rect 149716 50454 149744 70366
rect 149808 51814 149836 71402
rect 149900 53106 149928 71606
rect 150176 66910 150204 75618
rect 150452 73001 150480 79698
rect 150544 73154 150572 79784
rect 150866 79744 150894 80036
rect 150636 79716 150894 79744
rect 150636 78169 150664 79716
rect 150958 79642 150986 80036
rect 151050 79966 151078 80036
rect 151142 79966 151170 80036
rect 151038 79960 151090 79966
rect 151038 79902 151090 79908
rect 151130 79960 151182 79966
rect 151234 79937 151262 80036
rect 151326 79966 151354 80036
rect 151418 79966 151446 80036
rect 151510 79971 151538 80036
rect 151314 79960 151366 79966
rect 151130 79902 151182 79908
rect 151220 79928 151276 79937
rect 151314 79902 151366 79908
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151496 79962 151552 79971
rect 151602 79966 151630 80036
rect 151496 79897 151552 79906
rect 151590 79960 151642 79966
rect 151590 79902 151642 79908
rect 151220 79863 151276 79872
rect 151268 79824 151320 79830
rect 151694 79812 151722 80036
rect 151268 79766 151320 79772
rect 151648 79784 151722 79812
rect 150808 79620 150860 79626
rect 150808 79562 150860 79568
rect 150912 79614 150986 79642
rect 151084 79620 151136 79626
rect 150716 79552 150768 79558
rect 150716 79494 150768 79500
rect 150622 78160 150678 78169
rect 150622 78095 150678 78104
rect 150544 73126 150664 73154
rect 150438 72992 150494 73001
rect 150438 72927 150494 72936
rect 150636 69465 150664 73126
rect 150728 70038 150756 79494
rect 150820 72962 150848 79562
rect 150912 74089 150940 79614
rect 151084 79562 151136 79568
rect 151096 76022 151124 79562
rect 151176 79416 151228 79422
rect 151176 79358 151228 79364
rect 151188 79150 151216 79358
rect 151176 79144 151228 79150
rect 151176 79086 151228 79092
rect 151174 78296 151230 78305
rect 151174 78231 151230 78240
rect 151084 76016 151136 76022
rect 151084 75958 151136 75964
rect 151084 75880 151136 75886
rect 151084 75822 151136 75828
rect 150898 74080 150954 74089
rect 150898 74015 150954 74024
rect 150808 72956 150860 72962
rect 150808 72898 150860 72904
rect 151096 71534 151124 75822
rect 151084 71528 151136 71534
rect 151084 71470 151136 71476
rect 150716 70032 150768 70038
rect 150716 69974 150768 69980
rect 150622 69456 150678 69465
rect 150622 69391 150678 69400
rect 150164 66904 150216 66910
rect 150164 66846 150216 66852
rect 149888 53100 149940 53106
rect 149888 53042 149940 53048
rect 149796 51808 149848 51814
rect 149796 51750 149848 51756
rect 149704 50448 149756 50454
rect 149704 50390 149756 50396
rect 148324 40724 148376 40730
rect 148324 40666 148376 40672
rect 147772 28960 147824 28966
rect 147772 28902 147824 28908
rect 151096 14550 151124 71470
rect 151188 64705 151216 78231
rect 151280 65618 151308 79766
rect 151544 79688 151596 79694
rect 151648 79665 151676 79784
rect 151786 79744 151814 80036
rect 151878 79971 151906 80036
rect 151864 79962 151920 79971
rect 151864 79897 151920 79906
rect 151970 79898 151998 80036
rect 152062 79898 152090 80036
rect 152154 79971 152182 80036
rect 152140 79962 152196 79971
rect 151958 79892 152010 79898
rect 151958 79834 152010 79840
rect 152050 79892 152102 79898
rect 152140 79897 152196 79906
rect 152246 79898 152274 80036
rect 152338 79971 152366 80036
rect 152324 79962 152380 79971
rect 152430 79966 152458 80036
rect 152050 79834 152102 79840
rect 152234 79892 152286 79898
rect 152324 79897 152380 79906
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152234 79834 152286 79840
rect 152522 79801 152550 80036
rect 152614 79937 152642 80036
rect 152600 79928 152656 79937
rect 152706 79898 152734 80036
rect 152798 79966 152826 80036
rect 152890 79966 152918 80036
rect 152786 79960 152838 79966
rect 152786 79902 152838 79908
rect 152878 79960 152930 79966
rect 152878 79902 152930 79908
rect 152982 79898 153010 80036
rect 153074 79937 153102 80036
rect 153166 79966 153194 80036
rect 153154 79960 153206 79966
rect 153060 79928 153116 79937
rect 152600 79863 152656 79872
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 152970 79892 153022 79898
rect 153154 79902 153206 79908
rect 153258 79898 153286 80036
rect 153350 79971 153378 80036
rect 153336 79962 153392 79971
rect 153442 79966 153470 80036
rect 153534 79971 153562 80036
rect 153060 79863 153116 79872
rect 153246 79892 153298 79898
rect 153336 79897 153392 79906
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153520 79962 153576 79971
rect 153520 79897 153576 79906
rect 152970 79834 153022 79840
rect 153246 79834 153298 79840
rect 152370 79792 152426 79801
rect 151740 79716 151814 79744
rect 152188 79756 152240 79762
rect 151544 79630 151596 79636
rect 151634 79656 151690 79665
rect 151358 79520 151414 79529
rect 151358 79455 151414 79464
rect 151372 76106 151400 79455
rect 151556 77625 151584 79630
rect 151634 79591 151690 79600
rect 151636 79552 151688 79558
rect 151636 79494 151688 79500
rect 151542 77616 151598 77625
rect 151542 77551 151598 77560
rect 151372 76078 151492 76106
rect 151360 76016 151412 76022
rect 151360 75958 151412 75964
rect 151372 70174 151400 75958
rect 151464 74050 151492 76078
rect 151648 75886 151676 79494
rect 151740 77761 151768 79716
rect 152370 79727 152426 79736
rect 152508 79792 152564 79801
rect 152508 79727 152564 79736
rect 152648 79756 152700 79762
rect 152188 79698 152240 79704
rect 151910 79656 151966 79665
rect 151966 79614 152044 79642
rect 151910 79591 151966 79600
rect 151820 79552 151872 79558
rect 151820 79494 151872 79500
rect 151726 77752 151782 77761
rect 151726 77687 151782 77696
rect 151636 75880 151688 75886
rect 151636 75822 151688 75828
rect 151452 74044 151504 74050
rect 151452 73986 151504 73992
rect 151832 72554 151860 79494
rect 151912 79416 151964 79422
rect 151912 79358 151964 79364
rect 151924 72894 151952 79358
rect 151912 72888 151964 72894
rect 151912 72830 151964 72836
rect 151820 72548 151872 72554
rect 151820 72490 151872 72496
rect 151832 70394 151860 72490
rect 151832 70366 151952 70394
rect 151360 70168 151412 70174
rect 151360 70110 151412 70116
rect 151268 65612 151320 65618
rect 151268 65554 151320 65560
rect 151174 64696 151230 64705
rect 151174 64631 151230 64640
rect 151084 14544 151136 14550
rect 151084 14486 151136 14492
rect 151924 4690 151952 70366
rect 152016 70106 152044 79614
rect 152200 76650 152228 79698
rect 152278 79656 152334 79665
rect 152278 79591 152334 79600
rect 152108 76622 152228 76650
rect 152108 73166 152136 76622
rect 152096 73160 152148 73166
rect 152292 73154 152320 79591
rect 152384 74186 152412 79727
rect 152648 79698 152700 79704
rect 153016 79756 153068 79762
rect 153016 79698 153068 79704
rect 153476 79756 153528 79762
rect 153626 79744 153654 80036
rect 153718 79971 153746 80036
rect 153704 79962 153760 79971
rect 153704 79897 153760 79906
rect 153810 79898 153838 80036
rect 153902 79971 153930 80036
rect 153888 79962 153944 79971
rect 153798 79892 153850 79898
rect 153888 79897 153944 79906
rect 153994 79898 154022 80036
rect 154086 79937 154114 80036
rect 154178 79966 154206 80036
rect 154270 79966 154298 80036
rect 154166 79960 154218 79966
rect 154072 79928 154128 79937
rect 153798 79834 153850 79840
rect 153982 79892 154034 79898
rect 154166 79902 154218 79908
rect 154258 79960 154310 79966
rect 154258 79902 154310 79908
rect 154072 79863 154128 79872
rect 153982 79834 154034 79840
rect 153936 79756 153988 79762
rect 153626 79716 153700 79744
rect 153476 79698 153528 79704
rect 152554 79656 152610 79665
rect 152554 79591 152610 79600
rect 152660 79608 152688 79698
rect 152832 79688 152884 79694
rect 152832 79630 152884 79636
rect 152924 79688 152976 79694
rect 152924 79630 152976 79636
rect 152464 79348 152516 79354
rect 152464 79290 152516 79296
rect 152476 78334 152504 79290
rect 152464 78328 152516 78334
rect 152464 78270 152516 78276
rect 152372 74180 152424 74186
rect 152372 74122 152424 74128
rect 152096 73102 152148 73108
rect 152200 73126 152320 73154
rect 152200 70145 152228 73126
rect 152462 71768 152518 71777
rect 152462 71703 152518 71712
rect 152186 70136 152242 70145
rect 152004 70100 152056 70106
rect 152186 70071 152242 70080
rect 152004 70042 152056 70048
rect 152476 8294 152504 71703
rect 152568 68270 152596 79591
rect 152660 79580 152780 79608
rect 152648 79484 152700 79490
rect 152648 79426 152700 79432
rect 152660 71777 152688 79426
rect 152646 71768 152702 71777
rect 152646 71703 152702 71712
rect 152752 69018 152780 79580
rect 152844 75818 152872 79630
rect 152936 77178 152964 79630
rect 153028 79082 153056 79698
rect 153108 79688 153160 79694
rect 153108 79630 153160 79636
rect 153384 79688 153436 79694
rect 153384 79630 153436 79636
rect 153016 79076 153068 79082
rect 153016 79018 153068 79024
rect 152924 77172 152976 77178
rect 152924 77114 152976 77120
rect 152832 75812 152884 75818
rect 152832 75754 152884 75760
rect 153120 73681 153148 79630
rect 153396 78248 153424 79630
rect 153488 78316 153516 79698
rect 153488 78288 153608 78316
rect 153396 78220 153516 78248
rect 153384 78124 153436 78130
rect 153384 78066 153436 78072
rect 153290 78024 153346 78033
rect 153290 77959 153346 77968
rect 153106 73672 153162 73681
rect 153106 73607 153162 73616
rect 153304 72826 153332 77959
rect 153292 72820 153344 72826
rect 153292 72762 153344 72768
rect 152740 69012 152792 69018
rect 152740 68954 152792 68960
rect 152556 68264 152608 68270
rect 152556 68206 152608 68212
rect 153396 66026 153424 78066
rect 153488 69465 153516 78220
rect 153580 75041 153608 78288
rect 153672 78010 153700 79716
rect 153936 79698 153988 79704
rect 154120 79756 154172 79762
rect 154362 79744 154390 80036
rect 154454 79971 154482 80036
rect 154440 79962 154496 79971
rect 154440 79897 154496 79906
rect 154546 79812 154574 80036
rect 154638 79966 154666 80036
rect 154730 79971 154758 80036
rect 154626 79960 154678 79966
rect 154626 79902 154678 79908
rect 154716 79962 154772 79971
rect 154716 79897 154772 79906
rect 154822 79898 154850 80036
rect 154914 79966 154942 80036
rect 155006 79966 155034 80036
rect 155098 79966 155126 80036
rect 155190 79971 155218 80036
rect 154902 79960 154954 79966
rect 154902 79902 154954 79908
rect 154994 79960 155046 79966
rect 154994 79902 155046 79908
rect 155086 79960 155138 79966
rect 155086 79902 155138 79908
rect 155176 79962 155232 79971
rect 155282 79966 155310 80036
rect 155374 79966 155402 80036
rect 154810 79892 154862 79898
rect 155176 79897 155232 79906
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 155362 79960 155414 79966
rect 155362 79902 155414 79908
rect 154810 79834 154862 79840
rect 155466 79830 155494 80036
rect 155558 79971 155586 80036
rect 155544 79962 155600 79971
rect 155650 79966 155678 80036
rect 155742 79966 155770 80036
rect 155834 79966 155862 80036
rect 155926 79966 155954 80036
rect 156018 79966 156046 80036
rect 156110 79966 156138 80036
rect 156202 79966 156230 80036
rect 155544 79897 155600 79906
rect 155638 79960 155690 79966
rect 155638 79902 155690 79908
rect 155730 79960 155782 79966
rect 155730 79902 155782 79908
rect 155822 79960 155874 79966
rect 155822 79902 155874 79908
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 156006 79960 156058 79966
rect 156006 79902 156058 79908
rect 156098 79960 156150 79966
rect 156098 79902 156150 79908
rect 156190 79960 156242 79966
rect 156190 79902 156242 79908
rect 154120 79698 154172 79704
rect 154224 79716 154390 79744
rect 154500 79784 154574 79812
rect 155454 79824 155506 79830
rect 153752 79688 153804 79694
rect 153752 79630 153804 79636
rect 153764 78985 153792 79630
rect 153948 79490 153976 79698
rect 154026 79656 154082 79665
rect 154026 79591 154082 79600
rect 153936 79484 153988 79490
rect 153936 79426 153988 79432
rect 153750 78976 153806 78985
rect 153750 78911 153806 78920
rect 154040 78010 154068 79591
rect 154132 78130 154160 79698
rect 154120 78124 154172 78130
rect 154120 78066 154172 78072
rect 153672 77982 153884 78010
rect 154040 77982 154160 78010
rect 153752 76628 153804 76634
rect 153752 76570 153804 76576
rect 153566 75032 153622 75041
rect 153566 74967 153622 74976
rect 153474 69456 153530 69465
rect 153474 69391 153530 69400
rect 153384 66020 153436 66026
rect 153384 65962 153436 65968
rect 153764 64734 153792 76570
rect 153856 72350 153884 77982
rect 154028 77920 154080 77926
rect 154028 77862 154080 77868
rect 153936 74656 153988 74662
rect 153936 74598 153988 74604
rect 153844 72344 153896 72350
rect 153844 72286 153896 72292
rect 153948 72162 153976 74598
rect 153856 72134 153976 72162
rect 153856 71602 153884 72134
rect 153936 72072 153988 72078
rect 153936 72014 153988 72020
rect 153844 71596 153896 71602
rect 153844 71538 153896 71544
rect 153752 64728 153804 64734
rect 153752 64670 153804 64676
rect 153856 17270 153884 71538
rect 153948 65822 153976 72014
rect 153936 65816 153988 65822
rect 153936 65758 153988 65764
rect 154040 63510 154068 77862
rect 154132 64394 154160 77982
rect 154224 74662 154252 79716
rect 154304 79416 154356 79422
rect 154304 79358 154356 79364
rect 154316 75954 154344 79358
rect 154500 76634 154528 79784
rect 155454 79766 155506 79772
rect 155592 79824 155644 79830
rect 155592 79766 155644 79772
rect 155914 79824 155966 79830
rect 155966 79784 156046 79812
rect 155914 79766 155966 79772
rect 156018 79778 156046 79784
rect 156294 79778 156322 80036
rect 156386 79966 156414 80036
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156478 79830 156506 80036
rect 154856 79756 154908 79762
rect 154856 79698 154908 79704
rect 154580 79688 154632 79694
rect 154764 79688 154816 79694
rect 154580 79630 154632 79636
rect 154762 79656 154764 79665
rect 154816 79656 154818 79665
rect 154592 78674 154620 79630
rect 154672 79620 154724 79626
rect 154762 79591 154818 79600
rect 154672 79562 154724 79568
rect 154580 78668 154632 78674
rect 154580 78610 154632 78616
rect 154684 77217 154712 79562
rect 154762 79520 154818 79529
rect 154762 79455 154818 79464
rect 154670 77208 154726 77217
rect 154670 77143 154726 77152
rect 154488 76628 154540 76634
rect 154488 76570 154540 76576
rect 154672 76628 154724 76634
rect 154672 76570 154724 76576
rect 154304 75948 154356 75954
rect 154304 75890 154356 75896
rect 154212 74656 154264 74662
rect 154212 74598 154264 74604
rect 154316 73154 154344 75890
rect 154224 73126 154344 73154
rect 154224 72078 154252 73126
rect 154212 72072 154264 72078
rect 154212 72014 154264 72020
rect 154684 70310 154712 76570
rect 154776 73154 154804 79455
rect 154868 76634 154896 79698
rect 155132 79688 155184 79694
rect 155132 79630 155184 79636
rect 155500 79688 155552 79694
rect 155500 79630 155552 79636
rect 154948 78668 155000 78674
rect 154948 78610 155000 78616
rect 154856 76628 154908 76634
rect 154856 76570 154908 76576
rect 154960 76158 154988 78610
rect 155144 76226 155172 79630
rect 155408 79620 155460 79626
rect 155408 79562 155460 79568
rect 155316 76492 155368 76498
rect 155316 76434 155368 76440
rect 155132 76220 155184 76226
rect 155132 76162 155184 76168
rect 154948 76152 155000 76158
rect 154948 76094 155000 76100
rect 154776 73126 154896 73154
rect 154672 70304 154724 70310
rect 154672 70246 154724 70252
rect 154120 64388 154172 64394
rect 154120 64330 154172 64336
rect 154028 63504 154080 63510
rect 154028 63446 154080 63452
rect 154132 45554 154160 64330
rect 154868 64190 154896 73126
rect 155328 68882 155356 76434
rect 155420 76401 155448 79562
rect 155406 76392 155462 76401
rect 155406 76327 155462 76336
rect 155408 76152 155460 76158
rect 155408 76094 155460 76100
rect 155316 68876 155368 68882
rect 155316 68818 155368 68824
rect 154856 64184 154908 64190
rect 154856 64126 154908 64132
rect 155420 56574 155448 76094
rect 155512 57866 155540 79630
rect 155604 78674 155632 79766
rect 155776 79756 155828 79762
rect 156018 79750 156092 79778
rect 155776 79698 155828 79704
rect 155684 79688 155736 79694
rect 155684 79630 155736 79636
rect 155592 78668 155644 78674
rect 155592 78610 155644 78616
rect 155696 78062 155724 79630
rect 155684 78056 155736 78062
rect 155684 77998 155736 78004
rect 155592 76220 155644 76226
rect 155592 76162 155644 76168
rect 155604 66094 155632 76162
rect 155788 75750 155816 79698
rect 155868 79688 155920 79694
rect 155868 79630 155920 79636
rect 155880 78470 155908 79630
rect 155960 79552 156012 79558
rect 155960 79494 156012 79500
rect 155868 78464 155920 78470
rect 155868 78406 155920 78412
rect 155972 76786 156000 79494
rect 156064 76974 156092 79750
rect 156144 79756 156196 79762
rect 156144 79698 156196 79704
rect 156248 79750 156322 79778
rect 156466 79824 156518 79830
rect 156466 79766 156518 79772
rect 156570 79778 156598 80036
rect 156662 79966 156690 80036
rect 156650 79960 156702 79966
rect 156650 79902 156702 79908
rect 156570 79750 156644 79778
rect 156052 76968 156104 76974
rect 156052 76910 156104 76916
rect 156156 76786 156184 79698
rect 155880 76758 156000 76786
rect 156064 76758 156184 76786
rect 155776 75744 155828 75750
rect 155776 75686 155828 75692
rect 155592 66088 155644 66094
rect 155592 66030 155644 66036
rect 155880 62014 155908 76758
rect 156064 76650 156092 76758
rect 156248 76650 156276 79750
rect 156328 79688 156380 79694
rect 156328 79630 156380 79636
rect 156512 79688 156564 79694
rect 156616 79676 156644 79750
rect 156754 79744 156782 80036
rect 156846 79812 156874 80036
rect 156938 79966 156966 80036
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 157030 79812 157058 80036
rect 156846 79784 156920 79812
rect 156754 79716 156828 79744
rect 156616 79648 156736 79676
rect 156512 79630 156564 79636
rect 155972 76622 156092 76650
rect 156156 76622 156276 76650
rect 155868 62008 155920 62014
rect 155868 61950 155920 61956
rect 155500 57860 155552 57866
rect 155500 57802 155552 57808
rect 155408 56568 155460 56574
rect 155408 56510 155460 56516
rect 153948 45526 154160 45554
rect 153948 35222 153976 45526
rect 153936 35216 153988 35222
rect 153936 35158 153988 35164
rect 155880 25566 155908 61950
rect 155972 37262 156000 76622
rect 156052 75472 156104 75478
rect 156052 75414 156104 75420
rect 156064 46918 156092 75414
rect 156156 48278 156184 76622
rect 156236 76152 156288 76158
rect 156236 76094 156288 76100
rect 156248 63374 156276 76094
rect 156340 66162 156368 79630
rect 156420 79620 156472 79626
rect 156420 79562 156472 79568
rect 156432 78713 156460 79562
rect 156418 78704 156474 78713
rect 156418 78639 156474 78648
rect 156524 77994 156552 79630
rect 156604 79552 156656 79558
rect 156604 79494 156656 79500
rect 156616 78577 156644 79494
rect 156602 78568 156658 78577
rect 156602 78503 156658 78512
rect 156604 78464 156656 78470
rect 156604 78406 156656 78412
rect 156512 77988 156564 77994
rect 156512 77930 156564 77936
rect 156420 76900 156472 76906
rect 156420 76842 156472 76848
rect 156432 76430 156460 76842
rect 156512 76628 156564 76634
rect 156512 76570 156564 76576
rect 156420 76424 156472 76430
rect 156420 76366 156472 76372
rect 156420 76220 156472 76226
rect 156420 76162 156472 76168
rect 156432 70922 156460 76162
rect 156524 72758 156552 76570
rect 156616 76226 156644 78406
rect 156604 76220 156656 76226
rect 156604 76162 156656 76168
rect 156602 73128 156658 73137
rect 156602 73063 156658 73072
rect 156512 72752 156564 72758
rect 156512 72694 156564 72700
rect 156510 71768 156566 71777
rect 156510 71703 156566 71712
rect 156524 71097 156552 71703
rect 156510 71088 156566 71097
rect 156510 71023 156566 71032
rect 156420 70916 156472 70922
rect 156420 70858 156472 70864
rect 156616 69562 156644 73063
rect 156708 71777 156736 79648
rect 156800 72962 156828 79716
rect 156892 79121 156920 79784
rect 156984 79784 157058 79812
rect 156878 79112 156934 79121
rect 156878 79047 156934 79056
rect 156880 77308 156932 77314
rect 156880 77250 156932 77256
rect 156788 72956 156840 72962
rect 156788 72898 156840 72904
rect 156788 72752 156840 72758
rect 156788 72694 156840 72700
rect 156694 71768 156750 71777
rect 156694 71703 156750 71712
rect 156800 71058 156828 72694
rect 156788 71052 156840 71058
rect 156788 70994 156840 71000
rect 156604 69556 156656 69562
rect 156604 69498 156656 69504
rect 156328 66156 156380 66162
rect 156328 66098 156380 66104
rect 156892 63442 156920 77250
rect 156984 76634 157012 79784
rect 157122 79744 157150 80036
rect 157214 79966 157242 80036
rect 157306 79966 157334 80036
rect 157202 79960 157254 79966
rect 157202 79902 157254 79908
rect 157294 79960 157346 79966
rect 157294 79902 157346 79908
rect 157076 79716 157150 79744
rect 157248 79756 157300 79762
rect 156972 76628 157024 76634
rect 156972 76570 157024 76576
rect 157076 75478 157104 79716
rect 157248 79698 157300 79704
rect 157154 79656 157210 79665
rect 157154 79591 157210 79600
rect 157064 75472 157116 75478
rect 157064 75414 157116 75420
rect 157168 75002 157196 79591
rect 157260 78198 157288 79698
rect 157398 79676 157426 80036
rect 157490 79898 157518 80036
rect 157582 79937 157610 80036
rect 157568 79928 157624 79937
rect 157478 79892 157530 79898
rect 157568 79863 157624 79872
rect 157478 79834 157530 79840
rect 157674 79778 157702 80036
rect 157766 79812 157794 80036
rect 157858 79971 157886 80036
rect 157844 79962 157900 79971
rect 157844 79897 157900 79906
rect 157950 79898 157978 80036
rect 157938 79892 157990 79898
rect 157938 79834 157990 79840
rect 157766 79784 157840 79812
rect 157628 79762 157702 79778
rect 157616 79756 157702 79762
rect 157668 79750 157702 79756
rect 157616 79698 157668 79704
rect 157398 79648 157564 79676
rect 157340 79484 157392 79490
rect 157340 79426 157392 79432
rect 157248 78192 157300 78198
rect 157248 78134 157300 78140
rect 157352 76158 157380 79426
rect 157432 79348 157484 79354
rect 157432 79290 157484 79296
rect 157340 76152 157392 76158
rect 157340 76094 157392 76100
rect 157156 74996 157208 75002
rect 157156 74938 157208 74944
rect 157444 66745 157472 79290
rect 157536 68746 157564 79648
rect 157616 79620 157668 79626
rect 157616 79562 157668 79568
rect 157628 72282 157656 79562
rect 157708 79552 157760 79558
rect 157708 79494 157760 79500
rect 157720 77790 157748 79494
rect 157708 77784 157760 77790
rect 157708 77726 157760 77732
rect 157708 76968 157760 76974
rect 157708 76910 157760 76916
rect 157616 72276 157668 72282
rect 157616 72218 157668 72224
rect 157524 68740 157576 68746
rect 157524 68682 157576 68688
rect 157430 66736 157486 66745
rect 157430 66671 157486 66680
rect 157720 63986 157748 76910
rect 157812 73154 157840 79784
rect 157890 79792 157946 79801
rect 158042 79778 158070 80036
rect 158134 79966 158162 80036
rect 158226 79971 158254 80036
rect 158122 79960 158174 79966
rect 158122 79902 158174 79908
rect 158212 79962 158268 79971
rect 158212 79897 158268 79906
rect 158168 79824 158220 79830
rect 158166 79792 158168 79801
rect 158318 79812 158346 80036
rect 158220 79792 158222 79801
rect 158042 79750 158116 79778
rect 157890 79727 157946 79736
rect 157904 78062 157932 79727
rect 157984 79688 158036 79694
rect 157984 79630 158036 79636
rect 157996 78305 158024 79630
rect 157982 78296 158038 78305
rect 157982 78231 158038 78240
rect 157892 78056 157944 78062
rect 157892 77998 157944 78004
rect 158088 76673 158116 79750
rect 158166 79727 158222 79736
rect 158272 79784 158346 79812
rect 158272 79608 158300 79784
rect 158410 79744 158438 80036
rect 158502 79966 158530 80036
rect 158594 79966 158622 80036
rect 158686 79966 158714 80036
rect 158490 79960 158542 79966
rect 158490 79902 158542 79908
rect 158582 79960 158634 79966
rect 158582 79902 158634 79908
rect 158674 79960 158726 79966
rect 158674 79902 158726 79908
rect 158778 79830 158806 80036
rect 158766 79824 158818 79830
rect 158870 79801 158898 80036
rect 158766 79766 158818 79772
rect 158856 79792 158912 79801
rect 158180 79580 158300 79608
rect 158364 79716 158438 79744
rect 158856 79727 158912 79736
rect 158180 78266 158208 79580
rect 158260 79484 158312 79490
rect 158260 79426 158312 79432
rect 158168 78260 158220 78266
rect 158168 78202 158220 78208
rect 158168 78124 158220 78130
rect 158168 78066 158220 78072
rect 158074 76664 158130 76673
rect 158074 76599 158130 76608
rect 158180 73166 158208 78066
rect 158272 76226 158300 79426
rect 158364 78878 158392 79716
rect 158812 79688 158864 79694
rect 158962 79676 158990 80036
rect 158812 79630 158864 79636
rect 158916 79648 158990 79676
rect 159054 79676 159082 80036
rect 159146 79744 159174 80036
rect 159238 79812 159266 80036
rect 159330 79966 159358 80036
rect 159422 79966 159450 80036
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159410 79960 159462 79966
rect 159410 79902 159462 79908
rect 159514 79812 159542 80036
rect 159606 79830 159634 80036
rect 159698 79966 159726 80036
rect 159686 79960 159738 79966
rect 159686 79902 159738 79908
rect 159238 79801 159312 79812
rect 159238 79792 159326 79801
rect 159238 79784 159270 79792
rect 159146 79716 159220 79744
rect 159468 79784 159542 79812
rect 159594 79824 159646 79830
rect 159270 79727 159326 79736
rect 159364 79756 159416 79762
rect 159054 79648 159128 79676
rect 158444 79620 158496 79626
rect 158444 79562 158496 79568
rect 158352 78872 158404 78878
rect 158352 78814 158404 78820
rect 158352 78668 158404 78674
rect 158352 78610 158404 78616
rect 158260 76220 158312 76226
rect 158260 76162 158312 76168
rect 158260 75540 158312 75546
rect 158260 75482 158312 75488
rect 158272 75070 158300 75482
rect 158260 75064 158312 75070
rect 158260 75006 158312 75012
rect 158168 73160 158220 73166
rect 157812 73126 158116 73154
rect 158088 65958 158116 73126
rect 158168 73102 158220 73108
rect 158364 72690 158392 78610
rect 158456 76673 158484 79562
rect 158536 79552 158588 79558
rect 158536 79494 158588 79500
rect 158442 76664 158498 76673
rect 158442 76599 158498 76608
rect 158548 76498 158576 79494
rect 158720 78872 158772 78878
rect 158720 78814 158772 78820
rect 158628 77240 158680 77246
rect 158628 77182 158680 77188
rect 158536 76492 158588 76498
rect 158536 76434 158588 76440
rect 158640 74390 158668 77182
rect 158732 76906 158760 78814
rect 158824 78130 158852 79630
rect 158916 79558 158944 79648
rect 158904 79552 158956 79558
rect 158904 79494 158956 79500
rect 158996 79552 159048 79558
rect 158996 79494 159048 79500
rect 158904 79416 158956 79422
rect 158904 79358 158956 79364
rect 158812 78124 158864 78130
rect 158812 78066 158864 78072
rect 158720 76900 158772 76906
rect 158720 76842 158772 76848
rect 158720 76220 158772 76226
rect 158720 76162 158772 76168
rect 158628 74384 158680 74390
rect 158628 74326 158680 74332
rect 158628 73160 158680 73166
rect 158628 73102 158680 73108
rect 158352 72684 158404 72690
rect 158352 72626 158404 72632
rect 158364 70394 158392 72626
rect 158640 72418 158668 73102
rect 158628 72412 158680 72418
rect 158628 72354 158680 72360
rect 158364 70366 158576 70394
rect 158444 68060 158496 68066
rect 158444 68002 158496 68008
rect 158076 65952 158128 65958
rect 158076 65894 158128 65900
rect 158456 64870 158484 68002
rect 158444 64864 158496 64870
rect 158444 64806 158496 64812
rect 157708 63980 157760 63986
rect 157708 63922 157760 63928
rect 156880 63436 156932 63442
rect 156880 63378 156932 63384
rect 156236 63368 156288 63374
rect 156236 63310 156288 63316
rect 156144 48272 156196 48278
rect 156144 48214 156196 48220
rect 156052 46912 156104 46918
rect 156052 46854 156104 46860
rect 155960 37256 156012 37262
rect 155960 37198 156012 37204
rect 158548 33114 158576 70366
rect 158536 33108 158588 33114
rect 158536 33050 158588 33056
rect 155868 25560 155920 25566
rect 155868 25502 155920 25508
rect 153844 17264 153896 17270
rect 153844 17206 153896 17212
rect 152464 8288 152516 8294
rect 152464 8230 152516 8236
rect 152648 4888 152700 4894
rect 152648 4830 152700 4836
rect 148784 4684 148836 4690
rect 148784 4626 148836 4632
rect 151912 4684 151964 4690
rect 151912 4626 151964 4632
rect 146944 3528 146996 3534
rect 146944 3470 146996 3476
rect 148796 480 148824 4626
rect 152660 480 152688 4830
rect 158640 4826 158668 72354
rect 158732 62082 158760 76162
rect 158810 75984 158866 75993
rect 158810 75919 158866 75928
rect 158824 64841 158852 75919
rect 158916 66230 158944 79358
rect 159008 76090 159036 79494
rect 159100 76752 159128 79648
rect 159192 76820 159220 79716
rect 159364 79698 159416 79704
rect 159270 79656 159326 79665
rect 159270 79591 159326 79600
rect 159284 77110 159312 79591
rect 159272 77104 159324 77110
rect 159272 77046 159324 77052
rect 159192 76792 159312 76820
rect 159100 76724 159220 76752
rect 159088 76220 159140 76226
rect 159088 76162 159140 76168
rect 158996 76084 159048 76090
rect 158996 76026 159048 76032
rect 158996 75948 159048 75954
rect 158996 75890 159048 75896
rect 158904 66224 158956 66230
rect 158904 66166 158956 66172
rect 159008 65521 159036 75890
rect 159100 67658 159128 76162
rect 159192 68406 159220 76724
rect 159284 75954 159312 76792
rect 159376 76226 159404 79698
rect 159468 77314 159496 79784
rect 159594 79766 159646 79772
rect 159548 79688 159600 79694
rect 159790 79676 159818 80036
rect 159882 79966 159910 80036
rect 159974 79966 160002 80036
rect 160066 79966 160094 80036
rect 159870 79960 159922 79966
rect 159870 79902 159922 79908
rect 159962 79960 160014 79966
rect 159962 79902 160014 79908
rect 160054 79960 160106 79966
rect 160054 79902 160106 79908
rect 160158 79812 160186 80036
rect 159548 79630 159600 79636
rect 159744 79648 159818 79676
rect 159928 79784 160186 79812
rect 159456 77308 159508 77314
rect 159456 77250 159508 77256
rect 159456 77104 159508 77110
rect 159456 77046 159508 77052
rect 159364 76220 159416 76226
rect 159364 76162 159416 76168
rect 159364 76084 159416 76090
rect 159364 76026 159416 76032
rect 159272 75948 159324 75954
rect 159272 75890 159324 75896
rect 159376 68921 159404 76026
rect 159468 74322 159496 77046
rect 159456 74316 159508 74322
rect 159456 74258 159508 74264
rect 159560 71774 159588 79630
rect 159640 79620 159692 79626
rect 159640 79562 159692 79568
rect 159652 79393 159680 79562
rect 159638 79384 159694 79393
rect 159638 79319 159694 79328
rect 159744 74050 159772 79648
rect 159824 79552 159876 79558
rect 159824 79494 159876 79500
rect 159836 77081 159864 79494
rect 159822 77072 159878 77081
rect 159822 77007 159878 77016
rect 159928 75954 159956 79784
rect 160250 79744 160278 80036
rect 160342 79966 160370 80036
rect 160434 79966 160462 80036
rect 160526 79966 160554 80036
rect 160618 79966 160646 80036
rect 160710 79966 160738 80036
rect 160802 79966 160830 80036
rect 160894 79966 160922 80036
rect 160330 79960 160382 79966
rect 160330 79902 160382 79908
rect 160422 79960 160474 79966
rect 160422 79902 160474 79908
rect 160514 79960 160566 79966
rect 160514 79902 160566 79908
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160698 79960 160750 79966
rect 160698 79902 160750 79908
rect 160790 79960 160842 79966
rect 160790 79902 160842 79908
rect 160882 79960 160934 79966
rect 160986 79937 161014 80036
rect 161078 79966 161106 80036
rect 161066 79960 161118 79966
rect 160882 79902 160934 79908
rect 160972 79928 161028 79937
rect 161170 79937 161198 80036
rect 161066 79902 161118 79908
rect 161156 79928 161212 79937
rect 160972 79863 161028 79872
rect 161156 79863 161212 79872
rect 160514 79824 160566 79830
rect 160566 79772 160600 79778
rect 160514 79766 160600 79772
rect 160526 79750 160600 79766
rect 160250 79716 160324 79744
rect 160192 79620 160244 79626
rect 160192 79562 160244 79568
rect 160008 79552 160060 79558
rect 160008 79494 160060 79500
rect 159916 75948 159968 75954
rect 159916 75890 159968 75896
rect 159732 74044 159784 74050
rect 159732 73986 159784 73992
rect 160020 73817 160048 79494
rect 160100 78668 160152 78674
rect 160100 78610 160152 78616
rect 160112 75857 160140 78610
rect 160098 75848 160154 75857
rect 160098 75783 160154 75792
rect 160006 73808 160062 73817
rect 160006 73743 160062 73752
rect 159560 71746 159772 71774
rect 159744 71641 159772 71746
rect 159730 71632 159786 71641
rect 159730 71567 159786 71576
rect 159362 68912 159418 68921
rect 159362 68847 159418 68856
rect 160008 68536 160060 68542
rect 160008 68478 160060 68484
rect 159180 68400 159232 68406
rect 159180 68342 159232 68348
rect 160020 67658 160048 68478
rect 159088 67652 159140 67658
rect 159088 67594 159140 67600
rect 160008 67652 160060 67658
rect 160008 67594 160060 67600
rect 158994 65512 159050 65521
rect 158994 65447 159050 65456
rect 158810 64832 158866 64841
rect 158810 64767 158866 64776
rect 158720 62076 158772 62082
rect 158720 62018 158772 62024
rect 160020 18698 160048 67594
rect 160204 65346 160232 79562
rect 160296 78674 160324 79716
rect 160468 79688 160520 79694
rect 160468 79630 160520 79636
rect 160374 79520 160430 79529
rect 160374 79455 160430 79464
rect 160284 78668 160336 78674
rect 160284 78610 160336 78616
rect 160388 78130 160416 79455
rect 160376 78124 160428 78130
rect 160376 78066 160428 78072
rect 160480 76106 160508 79630
rect 160572 77246 160600 79750
rect 161112 79756 161164 79762
rect 161262 79744 161290 80036
rect 161354 79812 161382 80036
rect 161446 79966 161474 80036
rect 161434 79960 161486 79966
rect 161434 79902 161486 79908
rect 161354 79784 161428 79812
rect 161538 79801 161566 80036
rect 161630 79966 161658 80036
rect 161722 79966 161750 80036
rect 161814 79966 161842 80036
rect 161618 79960 161670 79966
rect 161618 79902 161670 79908
rect 161710 79960 161762 79966
rect 161710 79902 161762 79908
rect 161802 79960 161854 79966
rect 161802 79902 161854 79908
rect 161906 79898 161934 80036
rect 161998 79966 162026 80036
rect 162090 79971 162118 80036
rect 161986 79960 162038 79966
rect 161986 79902 162038 79908
rect 162076 79962 162132 79971
rect 161894 79892 161946 79898
rect 162076 79897 162132 79906
rect 161894 79834 161946 79840
rect 161262 79716 161336 79744
rect 161112 79698 161164 79704
rect 160836 79688 160888 79694
rect 160836 79630 160888 79636
rect 160652 79620 160704 79626
rect 160652 79562 160704 79568
rect 160560 77240 160612 77246
rect 160560 77182 160612 77188
rect 160388 76078 160508 76106
rect 160284 75880 160336 75886
rect 160284 75822 160336 75828
rect 160296 67318 160324 75822
rect 160388 68134 160416 76078
rect 160466 75984 160522 75993
rect 160466 75919 160522 75928
rect 160560 75948 160612 75954
rect 160480 68950 160508 75919
rect 160560 75890 160612 75896
rect 160468 68944 160520 68950
rect 160468 68886 160520 68892
rect 160376 68128 160428 68134
rect 160376 68070 160428 68076
rect 160480 68066 160508 68886
rect 160468 68060 160520 68066
rect 160468 68002 160520 68008
rect 160572 67930 160600 75890
rect 160664 75546 160692 79562
rect 160848 75886 160876 79630
rect 161124 78713 161152 79698
rect 161204 79620 161256 79626
rect 161204 79562 161256 79568
rect 161110 78704 161166 78713
rect 161110 78639 161166 78648
rect 161216 78266 161244 79562
rect 161204 78260 161256 78266
rect 161204 78202 161256 78208
rect 160836 75880 160888 75886
rect 160836 75822 160888 75828
rect 160652 75540 160704 75546
rect 160652 75482 160704 75488
rect 161308 74866 161336 79716
rect 161296 74860 161348 74866
rect 161296 74802 161348 74808
rect 161400 71774 161428 79784
rect 161524 79792 161580 79801
rect 161938 79792 161994 79801
rect 161524 79727 161580 79736
rect 161756 79756 161808 79762
rect 161756 79698 161808 79704
rect 161848 79756 161900 79762
rect 162182 79778 162210 80036
rect 161938 79727 161994 79736
rect 162090 79750 162210 79778
rect 161848 79698 161900 79704
rect 161478 79656 161534 79665
rect 161478 79591 161534 79600
rect 161664 79620 161716 79626
rect 161492 79218 161520 79591
rect 161664 79562 161716 79568
rect 161572 79552 161624 79558
rect 161572 79494 161624 79500
rect 161480 79212 161532 79218
rect 161480 79154 161532 79160
rect 161584 71774 161612 79494
rect 161308 71746 161428 71774
rect 161492 71746 161612 71774
rect 161308 70394 161336 71746
rect 161216 70366 161336 70394
rect 160560 67924 160612 67930
rect 160560 67866 160612 67872
rect 160284 67312 160336 67318
rect 160284 67254 160336 67260
rect 160192 65340 160244 65346
rect 160192 65282 160244 65288
rect 161216 61946 161244 70366
rect 161388 68808 161440 68814
rect 161388 68750 161440 68756
rect 161296 68468 161348 68474
rect 161296 68410 161348 68416
rect 161308 67930 161336 68410
rect 161400 68134 161428 68750
rect 161388 68128 161440 68134
rect 161388 68070 161440 68076
rect 161296 67924 161348 67930
rect 161296 67866 161348 67872
rect 161204 61940 161256 61946
rect 161204 61882 161256 61888
rect 161216 61266 161244 61882
rect 160100 61260 160152 61266
rect 160100 61202 160152 61208
rect 161204 61260 161256 61266
rect 161204 61202 161256 61208
rect 160112 57254 160140 61202
rect 160100 57248 160152 57254
rect 160100 57190 160152 57196
rect 161308 42090 161336 67866
rect 161296 42084 161348 42090
rect 161296 42026 161348 42032
rect 161400 39370 161428 68070
rect 161492 63306 161520 71746
rect 161676 64462 161704 79562
rect 161768 76090 161796 79698
rect 161756 76084 161808 76090
rect 161756 76026 161808 76032
rect 161756 75948 161808 75954
rect 161756 75890 161808 75896
rect 161768 65686 161796 75890
rect 161860 67998 161888 79698
rect 161952 68678 161980 79727
rect 162090 79642 162118 79750
rect 162274 79642 162302 80036
rect 162366 79778 162394 80036
rect 162458 79966 162486 80036
rect 162550 79966 162578 80036
rect 162446 79960 162498 79966
rect 162446 79902 162498 79908
rect 162538 79960 162590 79966
rect 162538 79902 162590 79908
rect 162642 79778 162670 80036
rect 162734 79830 162762 80036
rect 162826 79966 162854 80036
rect 162918 79971 162946 80036
rect 162814 79960 162866 79966
rect 162814 79902 162866 79908
rect 162904 79962 162960 79971
rect 163010 79966 163038 80036
rect 163102 79966 163130 80036
rect 162904 79897 162960 79906
rect 162998 79960 163050 79966
rect 162998 79902 163050 79908
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 162366 79750 162440 79778
rect 162090 79614 162164 79642
rect 162274 79614 162348 79642
rect 162032 79552 162084 79558
rect 162032 79494 162084 79500
rect 162044 77217 162072 79494
rect 162030 77208 162086 77217
rect 162030 77143 162086 77152
rect 162136 75954 162164 79614
rect 162320 78334 162348 79614
rect 162308 78328 162360 78334
rect 162308 78270 162360 78276
rect 162124 75948 162176 75954
rect 162124 75890 162176 75896
rect 162320 74390 162348 78270
rect 162308 74384 162360 74390
rect 162308 74326 162360 74332
rect 162412 71774 162440 79750
rect 162492 79756 162544 79762
rect 162492 79698 162544 79704
rect 162596 79750 162670 79778
rect 162722 79824 162774 79830
rect 162722 79766 162774 79772
rect 163044 79824 163096 79830
rect 163194 79812 163222 80036
rect 163286 79966 163314 80036
rect 163274 79960 163326 79966
rect 163274 79902 163326 79908
rect 163044 79766 163096 79772
rect 163148 79784 163222 79812
rect 162320 71746 162440 71774
rect 161940 68672 161992 68678
rect 161940 68614 161992 68620
rect 162320 68202 162348 71746
rect 162308 68196 162360 68202
rect 162308 68138 162360 68144
rect 161848 67992 161900 67998
rect 161848 67934 161900 67940
rect 161756 65680 161808 65686
rect 161756 65622 161808 65628
rect 161664 64456 161716 64462
rect 161664 64398 161716 64404
rect 161480 63300 161532 63306
rect 161480 63242 161532 63248
rect 161860 60734 161888 67934
rect 162320 60734 162348 68138
rect 162504 63238 162532 79698
rect 162596 79529 162624 79750
rect 162676 79688 162728 79694
rect 162676 79630 162728 79636
rect 162950 79656 163006 79665
rect 162582 79520 162638 79529
rect 162582 79455 162638 79464
rect 162584 79416 162636 79422
rect 162584 79358 162636 79364
rect 162596 72894 162624 79358
rect 162688 78946 162716 79630
rect 162768 79620 162820 79626
rect 162950 79591 163006 79600
rect 162768 79562 162820 79568
rect 162676 78940 162728 78946
rect 162676 78882 162728 78888
rect 162674 78568 162730 78577
rect 162674 78503 162730 78512
rect 162688 73914 162716 78503
rect 162676 73908 162728 73914
rect 162676 73850 162728 73856
rect 162584 72888 162636 72894
rect 162584 72830 162636 72836
rect 162780 72826 162808 79562
rect 162768 72820 162820 72826
rect 162768 72762 162820 72768
rect 162768 68672 162820 68678
rect 162768 68614 162820 68620
rect 162780 68066 162808 68614
rect 162768 68060 162820 68066
rect 162768 68002 162820 68008
rect 162492 63232 162544 63238
rect 162492 63174 162544 63180
rect 161860 60706 162164 60734
rect 162320 60706 162716 60734
rect 162136 49706 162164 60706
rect 162124 49700 162176 49706
rect 162124 49642 162176 49648
rect 161388 39364 161440 39370
rect 161388 39306 161440 39312
rect 162688 29714 162716 60706
rect 162676 29708 162728 29714
rect 162676 29650 162728 29656
rect 160008 18692 160060 18698
rect 160008 18634 160060 18640
rect 160376 9104 160428 9110
rect 160376 9046 160428 9052
rect 158628 4820 158680 4826
rect 158628 4762 158680 4768
rect 160388 480 160416 9046
rect 162780 6186 162808 68002
rect 162860 64116 162912 64122
rect 162860 64058 162912 64064
rect 162872 62898 162900 64058
rect 162860 62892 162912 62898
rect 162860 62834 162912 62840
rect 162964 55214 162992 79591
rect 163056 64122 163084 79766
rect 163148 78334 163176 79784
rect 163378 79778 163406 80036
rect 163470 79971 163498 80036
rect 163456 79962 163512 79971
rect 163456 79897 163512 79906
rect 163332 79750 163406 79778
rect 163332 79676 163360 79750
rect 163562 79744 163590 80036
rect 163654 79966 163682 80036
rect 163642 79960 163694 79966
rect 163642 79902 163694 79908
rect 163746 79898 163774 80036
rect 163838 79966 163866 80036
rect 163826 79960 163878 79966
rect 163930 79937 163958 80036
rect 163826 79902 163878 79908
rect 163916 79928 163972 79937
rect 163734 79892 163786 79898
rect 163916 79863 163972 79872
rect 163734 79834 163786 79840
rect 163872 79824 163924 79830
rect 164022 79778 164050 80036
rect 164114 79966 164142 80036
rect 164102 79960 164154 79966
rect 164102 79902 164154 79908
rect 164206 79830 164234 80036
rect 164298 79937 164326 80036
rect 164284 79928 164340 79937
rect 164390 79898 164418 80036
rect 164482 79937 164510 80036
rect 164574 79966 164602 80036
rect 164666 79966 164694 80036
rect 164758 79966 164786 80036
rect 164562 79960 164614 79966
rect 164468 79928 164524 79937
rect 164284 79863 164340 79872
rect 164378 79892 164430 79898
rect 164562 79902 164614 79908
rect 164654 79960 164706 79966
rect 164654 79902 164706 79908
rect 164746 79960 164798 79966
rect 164746 79902 164798 79908
rect 164468 79863 164524 79872
rect 164378 79834 164430 79840
rect 163872 79766 163924 79772
rect 163516 79716 163590 79744
rect 163240 79648 163360 79676
rect 163412 79688 163464 79694
rect 163240 78402 163268 79648
rect 163412 79630 163464 79636
rect 163320 79552 163372 79558
rect 163320 79494 163372 79500
rect 163228 78396 163280 78402
rect 163228 78338 163280 78344
rect 163136 78328 163188 78334
rect 163136 78270 163188 78276
rect 163332 78010 163360 79494
rect 163148 77982 163360 78010
rect 163148 67561 163176 77982
rect 163228 77920 163280 77926
rect 163228 77862 163280 77868
rect 163134 67552 163190 67561
rect 163134 67487 163190 67496
rect 163240 67454 163268 77862
rect 163424 75138 163452 79630
rect 163516 76362 163544 79716
rect 163688 79688 163740 79694
rect 163688 79630 163740 79636
rect 163596 79620 163648 79626
rect 163596 79562 163648 79568
rect 163608 77654 163636 79562
rect 163596 77648 163648 77654
rect 163596 77590 163648 77596
rect 163504 76356 163556 76362
rect 163504 76298 163556 76304
rect 163412 75132 163464 75138
rect 163412 75074 163464 75080
rect 163228 67448 163280 67454
rect 163228 67390 163280 67396
rect 163700 67114 163728 79630
rect 163884 78441 163912 79766
rect 163976 79750 164050 79778
rect 164194 79824 164246 79830
rect 164850 79778 164878 80036
rect 164942 79966 164970 80036
rect 165034 79966 165062 80036
rect 165126 79971 165154 80036
rect 164930 79960 164982 79966
rect 164930 79902 164982 79908
rect 165022 79960 165074 79966
rect 165022 79902 165074 79908
rect 165112 79962 165168 79971
rect 165218 79966 165246 80036
rect 165310 79971 165338 80036
rect 165112 79897 165168 79906
rect 165206 79960 165258 79966
rect 165206 79902 165258 79908
rect 165296 79962 165352 79971
rect 165402 79966 165430 80036
rect 165296 79897 165352 79906
rect 165390 79960 165442 79966
rect 165494 79937 165522 80036
rect 165390 79902 165442 79908
rect 165480 79928 165536 79937
rect 165586 79898 165614 80036
rect 165678 79966 165706 80036
rect 165770 79966 165798 80036
rect 165862 79971 165890 80036
rect 165666 79960 165718 79966
rect 165666 79902 165718 79908
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165848 79962 165904 79971
rect 165480 79863 165536 79872
rect 165574 79892 165626 79898
rect 165848 79897 165904 79906
rect 165954 79898 165982 80036
rect 166046 79971 166074 80036
rect 166032 79962 166088 79971
rect 165574 79834 165626 79840
rect 165942 79892 165994 79898
rect 166032 79897 166088 79906
rect 165942 79834 165994 79840
rect 166138 79830 166166 80036
rect 165344 79824 165396 79830
rect 164194 79766 164246 79772
rect 164516 79756 164568 79762
rect 163870 78432 163926 78441
rect 163870 78367 163926 78376
rect 163976 77926 164004 79750
rect 164516 79698 164568 79704
rect 164804 79750 164878 79778
rect 165250 79792 165306 79801
rect 164976 79756 165028 79762
rect 164056 79688 164108 79694
rect 164240 79688 164292 79694
rect 164056 79630 164108 79636
rect 164146 79656 164202 79665
rect 163964 77920 164016 77926
rect 163964 77862 164016 77868
rect 163872 77308 163924 77314
rect 163872 77250 163924 77256
rect 163884 74118 163912 77250
rect 163872 74112 163924 74118
rect 163872 74054 163924 74060
rect 163688 67108 163740 67114
rect 163688 67050 163740 67056
rect 163044 64116 163096 64122
rect 163044 64058 163096 64064
rect 162952 55208 163004 55214
rect 162952 55150 163004 55156
rect 164068 51066 164096 79630
rect 164240 79630 164292 79636
rect 164146 79591 164202 79600
rect 164160 75914 164188 79591
rect 164252 79082 164280 79630
rect 164424 79620 164476 79626
rect 164424 79562 164476 79568
rect 164240 79076 164292 79082
rect 164240 79018 164292 79024
rect 164160 75886 164280 75914
rect 164252 75274 164280 75886
rect 164240 75268 164292 75274
rect 164240 75210 164292 75216
rect 164332 75200 164384 75206
rect 164332 75142 164384 75148
rect 164240 75064 164292 75070
rect 164240 75006 164292 75012
rect 164148 67108 164200 67114
rect 164148 67050 164200 67056
rect 164056 51060 164108 51066
rect 164056 51002 164108 51008
rect 164160 38010 164188 67050
rect 164252 52426 164280 75006
rect 164344 63102 164372 75142
rect 164436 66026 164464 79562
rect 164528 67250 164556 79698
rect 164608 79620 164660 79626
rect 164608 79562 164660 79568
rect 164620 78577 164648 79562
rect 164700 79552 164752 79558
rect 164700 79494 164752 79500
rect 164606 78568 164662 78577
rect 164606 78503 164662 78512
rect 164608 75268 164660 75274
rect 164608 75210 164660 75216
rect 164516 67244 164568 67250
rect 164516 67186 164568 67192
rect 164620 67182 164648 75210
rect 164712 73778 164740 79494
rect 164700 73772 164752 73778
rect 164700 73714 164752 73720
rect 164804 71058 164832 79750
rect 164976 79698 165028 79704
rect 165160 79756 165212 79762
rect 166126 79824 166178 79830
rect 165344 79766 165396 79772
rect 165710 79792 165766 79801
rect 165250 79727 165306 79736
rect 165160 79698 165212 79704
rect 164884 79688 164936 79694
rect 164884 79630 164936 79636
rect 164896 76537 164924 79630
rect 164988 76673 165016 79698
rect 165066 79656 165122 79665
rect 165066 79591 165122 79600
rect 165080 77518 165108 79591
rect 165068 77512 165120 77518
rect 165068 77454 165120 77460
rect 164974 76664 165030 76673
rect 164974 76599 165030 76608
rect 164882 76528 164938 76537
rect 164882 76463 164938 76472
rect 165172 75070 165200 79698
rect 165160 75064 165212 75070
rect 165160 75006 165212 75012
rect 165264 72865 165292 79727
rect 165356 75206 165384 79766
rect 165620 79756 165672 79762
rect 165986 79792 166042 79801
rect 165710 79727 165766 79736
rect 165804 79756 165856 79762
rect 165620 79698 165672 79704
rect 165632 79665 165660 79698
rect 165618 79656 165674 79665
rect 165436 79620 165488 79626
rect 165618 79591 165674 79600
rect 165436 79562 165488 79568
rect 165344 75200 165396 75206
rect 165344 75142 165396 75148
rect 165250 72856 165306 72865
rect 165250 72791 165306 72800
rect 165448 71466 165476 79562
rect 165620 79484 165672 79490
rect 165620 79426 165672 79432
rect 165528 78328 165580 78334
rect 165528 78270 165580 78276
rect 165540 76430 165568 78270
rect 165528 76424 165580 76430
rect 165528 76366 165580 76372
rect 165632 74186 165660 79426
rect 165724 76634 165752 79727
rect 166126 79766 166178 79772
rect 165986 79727 166042 79736
rect 165804 79698 165856 79704
rect 165816 78033 165844 79698
rect 165896 79688 165948 79694
rect 165896 79630 165948 79636
rect 165802 78024 165858 78033
rect 165802 77959 165858 77968
rect 165804 77716 165856 77722
rect 165804 77658 165856 77664
rect 165712 76628 165764 76634
rect 165712 76570 165764 76576
rect 165712 76492 165764 76498
rect 165712 76434 165764 76440
rect 165620 74180 165672 74186
rect 165620 74122 165672 74128
rect 165436 71460 165488 71466
rect 165436 71402 165488 71408
rect 164792 71052 164844 71058
rect 164792 70994 164844 71000
rect 165344 71052 165396 71058
rect 165344 70994 165396 71000
rect 165356 68377 165384 70994
rect 165342 68368 165398 68377
rect 165342 68303 165398 68312
rect 164608 67176 164660 67182
rect 164608 67118 164660 67124
rect 164424 66020 164476 66026
rect 164424 65962 164476 65968
rect 164332 63096 164384 63102
rect 164332 63038 164384 63044
rect 164240 52420 164292 52426
rect 164240 52362 164292 52368
rect 164148 38004 164200 38010
rect 164148 37946 164200 37952
rect 165356 35290 165384 68303
rect 165436 64048 165488 64054
rect 165436 63990 165488 63996
rect 165344 35284 165396 35290
rect 165344 35226 165396 35232
rect 165448 16590 165476 63990
rect 165528 63096 165580 63102
rect 165528 63038 165580 63044
rect 165436 16584 165488 16590
rect 165436 16526 165488 16532
rect 165540 7614 165568 63038
rect 165724 62966 165752 76434
rect 165816 64734 165844 77658
rect 165908 70310 165936 79630
rect 166000 78577 166028 79727
rect 166080 79688 166132 79694
rect 166230 79676 166258 80036
rect 166322 79830 166350 80036
rect 166414 79966 166442 80036
rect 166506 79966 166534 80036
rect 166598 79971 166626 80036
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166494 79960 166546 79966
rect 166494 79902 166546 79908
rect 166584 79962 166640 79971
rect 166690 79966 166718 80036
rect 166782 79966 166810 80036
rect 166584 79897 166640 79906
rect 166678 79960 166730 79966
rect 166678 79902 166730 79908
rect 166770 79960 166822 79966
rect 166770 79902 166822 79908
rect 166310 79824 166362 79830
rect 166874 79778 166902 80036
rect 166966 79801 166994 80036
rect 167058 79971 167086 80036
rect 167044 79962 167100 79971
rect 167150 79966 167178 80036
rect 167242 79966 167270 80036
rect 167044 79897 167100 79906
rect 167138 79960 167190 79966
rect 167138 79902 167190 79908
rect 167230 79960 167282 79966
rect 167230 79902 167282 79908
rect 167334 79898 167362 80036
rect 167426 79937 167454 80036
rect 167518 79966 167546 80036
rect 167506 79960 167558 79966
rect 167412 79928 167468 79937
rect 167322 79892 167374 79898
rect 167506 79902 167558 79908
rect 167610 79898 167638 80036
rect 167702 79966 167730 80036
rect 167794 79966 167822 80036
rect 167690 79960 167742 79966
rect 167690 79902 167742 79908
rect 167782 79960 167834 79966
rect 167886 79937 167914 80036
rect 167782 79902 167834 79908
rect 167872 79928 167928 79937
rect 167412 79863 167468 79872
rect 167598 79892 167650 79898
rect 167322 79834 167374 79840
rect 167872 79863 167928 79872
rect 167598 79834 167650 79840
rect 166310 79766 166362 79772
rect 166632 79756 166684 79762
rect 166632 79698 166684 79704
rect 166828 79750 166902 79778
rect 166952 79792 167008 79801
rect 166356 79688 166408 79694
rect 166230 79648 166304 79676
rect 166080 79630 166132 79636
rect 165986 78568 166042 78577
rect 165986 78503 166042 78512
rect 165988 78192 166040 78198
rect 165988 78134 166040 78140
rect 166000 73710 166028 78134
rect 165988 73704 166040 73710
rect 165988 73646 166040 73652
rect 165896 70304 165948 70310
rect 165896 70246 165948 70252
rect 166092 70174 166120 79630
rect 166172 78124 166224 78130
rect 166172 78066 166224 78072
rect 166184 71097 166212 78066
rect 166276 76226 166304 79648
rect 166356 79630 166408 79636
rect 166448 79688 166500 79694
rect 166448 79630 166500 79636
rect 166538 79656 166594 79665
rect 166368 77722 166396 79630
rect 166356 77716 166408 77722
rect 166356 77658 166408 77664
rect 166460 76294 166488 79630
rect 166538 79591 166540 79600
rect 166592 79591 166594 79600
rect 166540 79562 166592 79568
rect 166540 79416 166592 79422
rect 166540 79358 166592 79364
rect 166552 78470 166580 79358
rect 166644 78674 166672 79698
rect 166644 78646 166764 78674
rect 166540 78464 166592 78470
rect 166540 78406 166592 78412
rect 166552 77042 166580 78406
rect 166632 78396 166684 78402
rect 166632 78338 166684 78344
rect 166540 77036 166592 77042
rect 166540 76978 166592 76984
rect 166448 76288 166500 76294
rect 166448 76230 166500 76236
rect 166264 76220 166316 76226
rect 166264 76162 166316 76168
rect 166264 76084 166316 76090
rect 166264 76026 166316 76032
rect 166276 73030 166304 76026
rect 166644 74254 166672 78338
rect 166632 74248 166684 74254
rect 166632 74190 166684 74196
rect 166264 73024 166316 73030
rect 166264 72966 166316 72972
rect 166170 71088 166226 71097
rect 166170 71023 166226 71032
rect 166736 70394 166764 78646
rect 166828 76498 166856 79750
rect 166952 79727 167008 79736
rect 167276 79756 167328 79762
rect 167276 79698 167328 79704
rect 167000 79620 167052 79626
rect 167000 79562 167052 79568
rect 167184 79620 167236 79626
rect 167184 79562 167236 79568
rect 167012 78606 167040 79562
rect 167000 78600 167052 78606
rect 167000 78542 167052 78548
rect 166816 76492 166868 76498
rect 166816 76434 166868 76440
rect 166908 76220 166960 76226
rect 166908 76162 166960 76168
rect 166184 70366 166764 70394
rect 166080 70168 166132 70174
rect 166080 70110 166132 70116
rect 166092 69086 166120 70110
rect 166080 69080 166132 69086
rect 166080 69022 166132 69028
rect 165804 64728 165856 64734
rect 165804 64670 165856 64676
rect 165712 62960 165764 62966
rect 165712 62902 165764 62908
rect 166184 59294 166212 70366
rect 166264 69080 166316 69086
rect 166264 69022 166316 69028
rect 166172 59288 166224 59294
rect 166172 59230 166224 59236
rect 166276 58682 166304 69022
rect 166920 66978 166948 76162
rect 167196 75274 167224 79562
rect 167288 78266 167316 79698
rect 167460 79688 167512 79694
rect 167978 79676 168006 80036
rect 168070 79801 168098 80036
rect 168056 79792 168112 79801
rect 168056 79727 168112 79736
rect 168162 79744 168190 80036
rect 168254 79937 168282 80036
rect 168240 79928 168296 79937
rect 168240 79863 168296 79872
rect 168346 79812 168374 80036
rect 168438 79966 168466 80036
rect 168426 79960 168478 79966
rect 168426 79902 168478 79908
rect 168530 79898 168558 80036
rect 168622 79971 168650 80036
rect 168608 79962 168664 79971
rect 168518 79892 168570 79898
rect 168608 79897 168664 79906
rect 168518 79834 168570 79840
rect 168300 79784 168374 79812
rect 168162 79716 168236 79744
rect 167978 79648 168144 79676
rect 167460 79630 167512 79636
rect 167368 79620 167420 79626
rect 167368 79562 167420 79568
rect 167276 78260 167328 78266
rect 167276 78202 167328 78208
rect 167276 77920 167328 77926
rect 167276 77862 167328 77868
rect 167184 75268 167236 75274
rect 167184 75210 167236 75216
rect 167092 75200 167144 75206
rect 167092 75142 167144 75148
rect 166908 66972 166960 66978
rect 166908 66914 166960 66920
rect 167104 63034 167132 75142
rect 167184 74792 167236 74798
rect 167184 74734 167236 74740
rect 167196 65754 167224 74734
rect 167184 65748 167236 65754
rect 167184 65690 167236 65696
rect 167288 65618 167316 77862
rect 167380 67658 167408 79562
rect 167472 78130 167500 79630
rect 167552 79620 167604 79626
rect 167552 79562 167604 79568
rect 167828 79620 167880 79626
rect 167828 79562 167880 79568
rect 167460 78124 167512 78130
rect 167460 78066 167512 78072
rect 167564 77926 167592 79562
rect 167840 79064 167868 79562
rect 167920 79552 167972 79558
rect 167920 79494 167972 79500
rect 167656 79036 167868 79064
rect 167552 77920 167604 77926
rect 167552 77862 167604 77868
rect 167656 69630 167684 79036
rect 167826 78976 167882 78985
rect 167932 78946 167960 79494
rect 168116 79286 168144 79648
rect 168104 79280 168156 79286
rect 168104 79222 168156 79228
rect 167826 78911 167882 78920
rect 167920 78940 167972 78946
rect 167736 75268 167788 75274
rect 167736 75210 167788 75216
rect 167644 69624 167696 69630
rect 167644 69566 167696 69572
rect 167368 67652 167420 67658
rect 167368 67594 167420 67600
rect 167276 65612 167328 65618
rect 167276 65554 167328 65560
rect 167092 63028 167144 63034
rect 167092 62970 167144 62976
rect 166908 62960 166960 62966
rect 166908 62902 166960 62908
rect 166264 58676 166316 58682
rect 166264 58618 166316 58624
rect 166920 14482 166948 62902
rect 167104 60110 167132 62970
rect 167748 62762 167776 75210
rect 167840 69970 167868 78911
rect 167920 78882 167972 78888
rect 168208 78674 168236 79716
rect 168300 79422 168328 79784
rect 168714 79744 168742 80036
rect 168806 79966 168834 80036
rect 168898 79966 168926 80036
rect 168990 79966 169018 80036
rect 169082 79966 169110 80036
rect 168794 79960 168846 79966
rect 168794 79902 168846 79908
rect 168886 79960 168938 79966
rect 168886 79902 168938 79908
rect 168978 79960 169030 79966
rect 168978 79902 169030 79908
rect 169070 79960 169122 79966
rect 169070 79902 169122 79908
rect 168932 79824 168984 79830
rect 168932 79766 168984 79772
rect 168668 79716 168742 79744
rect 168840 79756 168892 79762
rect 168472 79688 168524 79694
rect 168472 79630 168524 79636
rect 168288 79416 168340 79422
rect 168288 79358 168340 79364
rect 168378 79248 168434 79257
rect 168378 79183 168434 79192
rect 168286 78976 168342 78985
rect 168286 78911 168342 78920
rect 168116 78646 168236 78674
rect 167920 77716 167972 77722
rect 167920 77658 167972 77664
rect 167828 69964 167880 69970
rect 167828 69906 167880 69912
rect 167932 63170 167960 77658
rect 168116 74798 168144 78646
rect 168196 78600 168248 78606
rect 168196 78542 168248 78548
rect 168104 74792 168156 74798
rect 168104 74734 168156 74740
rect 168104 68128 168156 68134
rect 168104 68070 168156 68076
rect 168116 67658 168144 68070
rect 168104 67652 168156 67658
rect 168104 67594 168156 67600
rect 167920 63164 167972 63170
rect 167920 63106 167972 63112
rect 167736 62756 167788 62762
rect 167736 62698 167788 62704
rect 168116 60734 168144 67594
rect 168208 67590 168236 78542
rect 168300 75206 168328 78911
rect 168392 78742 168420 79183
rect 168380 78736 168432 78742
rect 168380 78678 168432 78684
rect 168484 76702 168512 79630
rect 168564 79620 168616 79626
rect 168564 79562 168616 79568
rect 168576 78418 168604 79562
rect 168668 78674 168696 79716
rect 168840 79698 168892 79704
rect 168746 79656 168802 79665
rect 168746 79591 168802 79600
rect 168656 78668 168708 78674
rect 168656 78610 168708 78616
rect 168576 78390 168696 78418
rect 168564 78328 168616 78334
rect 168564 78270 168616 78276
rect 168472 76696 168524 76702
rect 168472 76638 168524 76644
rect 168472 75948 168524 75954
rect 168472 75890 168524 75896
rect 168288 75200 168340 75206
rect 168288 75142 168340 75148
rect 168196 67584 168248 67590
rect 168196 67526 168248 67532
rect 168288 65748 168340 65754
rect 168288 65690 168340 65696
rect 168116 60706 168236 60734
rect 167092 60104 167144 60110
rect 167092 60046 167144 60052
rect 168208 33794 168236 60706
rect 168196 33788 168248 33794
rect 168196 33730 168248 33736
rect 168300 31074 168328 65690
rect 168484 60722 168512 75890
rect 168576 62898 168604 78270
rect 168668 68649 168696 78390
rect 168760 75886 168788 79591
rect 168852 75954 168880 79698
rect 168840 75948 168892 75954
rect 168840 75890 168892 75896
rect 168748 75880 168800 75886
rect 168748 75822 168800 75828
rect 168654 68640 168710 68649
rect 168654 68575 168710 68584
rect 168944 68270 168972 79766
rect 169174 79676 169202 80036
rect 169266 79971 169294 80036
rect 169252 79962 169308 79971
rect 169358 79966 169386 80036
rect 169252 79897 169308 79906
rect 169346 79960 169398 79966
rect 169346 79902 169398 79908
rect 169450 79744 169478 80036
rect 169542 79812 169570 80036
rect 169634 79937 169662 80036
rect 169726 79966 169754 80036
rect 169714 79960 169766 79966
rect 169620 79928 169676 79937
rect 169714 79902 169766 79908
rect 169620 79863 169676 79872
rect 169668 79824 169720 79830
rect 169542 79784 169616 79812
rect 169450 79716 169524 79744
rect 169174 79648 169248 79676
rect 169024 79620 169076 79626
rect 169024 79562 169076 79568
rect 169036 77722 169064 79562
rect 169024 77716 169076 77722
rect 169024 77658 169076 77664
rect 169220 75410 169248 79648
rect 169392 79620 169444 79626
rect 169392 79562 169444 79568
rect 169300 78668 169352 78674
rect 169300 78610 169352 78616
rect 169312 78180 169340 78610
rect 169404 78334 169432 79562
rect 169496 78849 169524 79716
rect 169482 78840 169538 78849
rect 169482 78775 169538 78784
rect 169392 78328 169444 78334
rect 169392 78270 169444 78276
rect 169484 78192 169536 78198
rect 169312 78152 169432 78180
rect 169300 77988 169352 77994
rect 169300 77930 169352 77936
rect 169208 75404 169260 75410
rect 169208 75346 169260 75352
rect 169312 74526 169340 77930
rect 169300 74520 169352 74526
rect 169300 74462 169352 74468
rect 169404 71670 169432 78152
rect 169484 78134 169536 78140
rect 169496 72554 169524 78134
rect 169484 72548 169536 72554
rect 169484 72490 169536 72496
rect 169392 71664 169444 71670
rect 169392 71606 169444 71612
rect 169588 70394 169616 79784
rect 169818 79778 169846 80036
rect 169910 79966 169938 80036
rect 170002 79971 170030 80036
rect 169898 79960 169950 79966
rect 169898 79902 169950 79908
rect 169988 79962 170044 79971
rect 169988 79897 170044 79906
rect 170094 79778 170122 80036
rect 170186 79966 170214 80036
rect 170278 79971 170306 80036
rect 170174 79960 170226 79966
rect 170174 79902 170226 79908
rect 170264 79962 170320 79971
rect 170264 79897 170320 79906
rect 170370 79898 170398 80036
rect 170462 79966 170490 80036
rect 170554 79966 170582 80036
rect 170450 79960 170502 79966
rect 170450 79902 170502 79908
rect 170542 79960 170594 79966
rect 170542 79902 170594 79908
rect 170358 79892 170410 79898
rect 170358 79834 170410 79840
rect 170646 79812 170674 80036
rect 170738 79937 170766 80036
rect 170724 79928 170780 79937
rect 170724 79863 170780 79872
rect 170830 79812 170858 80036
rect 169668 79766 169720 79772
rect 169680 78334 169708 79766
rect 169772 79750 169846 79778
rect 169956 79750 170122 79778
rect 170600 79784 170674 79812
rect 170784 79784 170858 79812
rect 170312 79756 170364 79762
rect 169668 78328 169720 78334
rect 169668 78270 169720 78276
rect 169668 78056 169720 78062
rect 169668 77998 169720 78004
rect 169680 72457 169708 77998
rect 169772 76129 169800 79750
rect 169956 79744 169984 79750
rect 169910 79716 169984 79744
rect 169910 79676 169938 79716
rect 170312 79698 170364 79704
rect 170404 79756 170456 79762
rect 170404 79698 170456 79704
rect 169864 79648 169938 79676
rect 170036 79688 170088 79694
rect 169758 76120 169814 76129
rect 169758 76055 169814 76064
rect 169864 75914 169892 79648
rect 170036 79630 170088 79636
rect 170128 79688 170180 79694
rect 170128 79630 170180 79636
rect 170048 76294 170076 79630
rect 170036 76288 170088 76294
rect 170036 76230 170088 76236
rect 170034 75984 170090 75993
rect 169772 75886 169892 75914
rect 169944 75948 169996 75954
rect 170140 75954 170168 79630
rect 170324 77722 170352 79698
rect 170312 77716 170364 77722
rect 170312 77658 170364 77664
rect 170034 75919 170090 75928
rect 170128 75948 170180 75954
rect 169944 75890 169996 75896
rect 169666 72448 169722 72457
rect 169666 72383 169722 72392
rect 169588 70366 169708 70394
rect 168932 68264 168984 68270
rect 168932 68206 168984 68212
rect 168564 62892 168616 62898
rect 168564 62834 168616 62840
rect 168472 60716 168524 60722
rect 168472 60658 168524 60664
rect 169680 59362 169708 70366
rect 169668 59356 169720 59362
rect 169668 59298 169720 59304
rect 169772 57934 169800 75886
rect 169852 75812 169904 75818
rect 169852 75754 169904 75760
rect 169864 64870 169892 75754
rect 169852 64864 169904 64870
rect 169852 64806 169904 64812
rect 169956 64802 169984 75890
rect 170048 66094 170076 75919
rect 170128 75890 170180 75896
rect 170416 67046 170444 79698
rect 170496 79688 170548 79694
rect 170496 79630 170548 79636
rect 170508 78062 170536 79630
rect 170496 78056 170548 78062
rect 170496 77998 170548 78004
rect 170600 71774 170628 79784
rect 170680 79212 170732 79218
rect 170680 79154 170732 79160
rect 170692 76022 170720 79154
rect 170680 76016 170732 76022
rect 170680 75958 170732 75964
rect 170784 75614 170812 79784
rect 170922 79778 170950 80036
rect 171014 79898 171042 80036
rect 171106 79937 171134 80036
rect 171092 79928 171148 79937
rect 171002 79892 171054 79898
rect 171198 79898 171226 80036
rect 171290 79966 171318 80036
rect 171278 79960 171330 79966
rect 171278 79902 171330 79908
rect 171092 79863 171148 79872
rect 171186 79892 171238 79898
rect 171002 79834 171054 79840
rect 171186 79834 171238 79840
rect 171382 79812 171410 80036
rect 171138 79792 171194 79801
rect 170922 79750 171088 79778
rect 170956 79688 171008 79694
rect 170956 79630 171008 79636
rect 170862 78976 170918 78985
rect 170862 78911 170918 78920
rect 170876 75818 170904 78911
rect 170968 77926 170996 79630
rect 171060 79218 171088 79750
rect 171138 79727 171194 79736
rect 171336 79784 171410 79812
rect 171048 79212 171100 79218
rect 171048 79154 171100 79160
rect 171152 78878 171180 79727
rect 171230 79656 171286 79665
rect 171230 79591 171286 79600
rect 171244 79257 171272 79591
rect 171230 79248 171286 79257
rect 171230 79183 171286 79192
rect 171140 78872 171192 78878
rect 171140 78814 171192 78820
rect 170956 77920 171008 77926
rect 170956 77862 171008 77868
rect 170956 77648 171008 77654
rect 170956 77590 171008 77596
rect 170864 75812 170916 75818
rect 170864 75754 170916 75760
rect 170772 75608 170824 75614
rect 170772 75550 170824 75556
rect 170968 73137 170996 77590
rect 171336 77194 171364 79784
rect 171474 79744 171502 80036
rect 171566 79812 171594 80036
rect 171658 79966 171686 80036
rect 171646 79960 171698 79966
rect 171646 79902 171698 79908
rect 171566 79801 171640 79812
rect 171566 79792 171654 79801
rect 171566 79784 171598 79792
rect 171428 79716 171502 79744
rect 171750 79778 171778 80036
rect 171842 79898 171870 80036
rect 171934 79903 171962 80036
rect 171830 79892 171882 79898
rect 171830 79834 171882 79840
rect 171920 79894 171976 79903
rect 171920 79829 171976 79838
rect 172026 79812 172054 80036
rect 172118 79966 172146 80036
rect 172210 79966 172238 80036
rect 172302 79971 172330 80036
rect 172106 79960 172158 79966
rect 172106 79902 172158 79908
rect 172198 79960 172250 79966
rect 172198 79902 172250 79908
rect 172288 79962 172344 79971
rect 172394 79966 172422 80036
rect 172486 79971 172514 80036
rect 172288 79897 172344 79906
rect 172382 79960 172434 79966
rect 172382 79902 172434 79908
rect 172472 79962 172528 79971
rect 172578 79966 172606 80036
rect 172472 79897 172528 79906
rect 172566 79960 172618 79966
rect 172670 79937 172698 80036
rect 172566 79902 172618 79908
rect 172656 79928 172712 79937
rect 172656 79863 172712 79872
rect 172428 79824 172480 79830
rect 172026 79784 172100 79812
rect 171598 79727 171654 79736
rect 171704 79750 171778 79778
rect 171428 79506 171456 79716
rect 171600 79688 171652 79694
rect 171600 79630 171652 79636
rect 171428 79478 171548 79506
rect 171416 79416 171468 79422
rect 171416 79358 171468 79364
rect 171152 77166 171364 77194
rect 170954 73128 171010 73137
rect 170954 73063 171010 73072
rect 170508 71746 170628 71774
rect 170508 71534 170536 71746
rect 170496 71528 170548 71534
rect 170496 71470 170548 71476
rect 171152 68785 171180 77166
rect 171232 76084 171284 76090
rect 171232 76026 171284 76032
rect 171138 68776 171194 68785
rect 171138 68711 171194 68720
rect 170404 67040 170456 67046
rect 170404 66982 170456 66988
rect 170416 66366 170444 66982
rect 170404 66360 170456 66366
rect 170404 66302 170456 66308
rect 170956 66360 171008 66366
rect 170956 66302 171008 66308
rect 170036 66088 170088 66094
rect 170036 66030 170088 66036
rect 169944 64796 169996 64802
rect 169944 64738 169996 64744
rect 169760 57928 169812 57934
rect 169760 57870 169812 57876
rect 168288 31068 168340 31074
rect 168288 31010 168340 31016
rect 170968 28354 170996 66302
rect 171140 65612 171192 65618
rect 171140 65554 171192 65560
rect 171048 64864 171100 64870
rect 171048 64806 171100 64812
rect 171060 64394 171088 64806
rect 171048 64388 171100 64394
rect 171048 64330 171100 64336
rect 170956 28348 171008 28354
rect 170956 28290 171008 28296
rect 167000 26308 167052 26314
rect 167000 26250 167052 26256
rect 167012 16574 167040 26250
rect 171060 22846 171088 64330
rect 171048 22840 171100 22846
rect 171048 22782 171100 22788
rect 167012 16546 168144 16574
rect 166908 14476 166960 14482
rect 166908 14418 166960 14424
rect 165528 7608 165580 7614
rect 165528 7550 165580 7556
rect 162768 6180 162820 6186
rect 162768 6122 162820 6128
rect 168116 480 168144 16546
rect 110758 354 110870 480
rect 110432 326 110870 354
rect 99166 -960 99278 326
rect 103030 -960 103142 326
rect 106894 -960 107006 326
rect 110758 -960 110870 326
rect 113978 -960 114090 480
rect 117842 -960 117954 480
rect 121706 -960 121818 480
rect 125570 -960 125682 480
rect 129434 -960 129546 480
rect 133298 -960 133410 480
rect 137162 -960 137274 480
rect 141026 -960 141138 480
rect 144890 -960 145002 480
rect 148754 -960 148866 480
rect 152618 -960 152730 480
rect 156482 -960 156594 480
rect 160346 -960 160458 480
rect 164210 -960 164322 480
rect 168074 -960 168186 480
rect 171152 354 171180 65554
rect 171244 64870 171272 76026
rect 171324 75948 171376 75954
rect 171324 75890 171376 75896
rect 171336 69737 171364 75890
rect 171428 71602 171456 79358
rect 171416 71596 171468 71602
rect 171416 71538 171468 71544
rect 171520 71194 171548 79478
rect 171612 75818 171640 79630
rect 171704 75954 171732 79750
rect 171968 79688 172020 79694
rect 171968 79630 172020 79636
rect 171784 79620 171836 79626
rect 171784 79562 171836 79568
rect 171796 78470 171824 79562
rect 171784 78464 171836 78470
rect 171784 78406 171836 78412
rect 171980 77568 172008 79630
rect 172072 79490 172100 79784
rect 172612 79824 172664 79830
rect 172428 79766 172480 79772
rect 172518 79792 172574 79801
rect 172244 79756 172296 79762
rect 172244 79698 172296 79704
rect 172060 79484 172112 79490
rect 172060 79426 172112 79432
rect 172152 79212 172204 79218
rect 172152 79154 172204 79160
rect 172164 78996 172192 79154
rect 172072 78968 172192 78996
rect 172072 78742 172100 78968
rect 172060 78736 172112 78742
rect 172060 78678 172112 78684
rect 171888 77540 172008 77568
rect 171888 76090 171916 77540
rect 171876 76084 171928 76090
rect 171876 76026 171928 76032
rect 172060 76016 172112 76022
rect 171966 75984 172022 75993
rect 171692 75948 171744 75954
rect 172060 75958 172112 75964
rect 171966 75919 172022 75928
rect 171692 75890 171744 75896
rect 171784 75880 171836 75886
rect 171784 75822 171836 75828
rect 171600 75812 171652 75818
rect 171600 75754 171652 75760
rect 171796 71330 171824 75822
rect 171784 71324 171836 71330
rect 171784 71266 171836 71272
rect 171508 71188 171560 71194
rect 171508 71130 171560 71136
rect 171520 70394 171548 71130
rect 171520 70366 171824 70394
rect 171322 69728 171378 69737
rect 171322 69663 171378 69672
rect 171232 64864 171284 64870
rect 171232 64806 171284 64812
rect 171796 4894 171824 70366
rect 171980 69902 172008 75919
rect 172072 70106 172100 75958
rect 172256 75886 172284 79698
rect 172336 79688 172388 79694
rect 172336 79630 172388 79636
rect 172348 78810 172376 79630
rect 172336 78804 172388 78810
rect 172336 78746 172388 78752
rect 172440 77704 172468 79766
rect 172612 79766 172664 79772
rect 172518 79727 172574 79736
rect 172348 77676 172468 77704
rect 172244 75880 172296 75886
rect 172244 75822 172296 75828
rect 172348 73098 172376 77676
rect 172532 77602 172560 79727
rect 172440 77574 172560 77602
rect 172440 77110 172468 77574
rect 172520 77512 172572 77518
rect 172520 77454 172572 77460
rect 172428 77104 172480 77110
rect 172428 77046 172480 77052
rect 172532 73982 172560 77454
rect 172520 73976 172572 73982
rect 172520 73918 172572 73924
rect 172336 73092 172388 73098
rect 172336 73034 172388 73040
rect 172624 70378 172652 79766
rect 172762 79642 172790 80036
rect 172854 79744 172882 80036
rect 172946 79812 172974 80036
rect 173038 79966 173066 80036
rect 173130 79971 173158 80036
rect 173026 79960 173078 79966
rect 173026 79902 173078 79908
rect 173116 79962 173172 79971
rect 173116 79897 173172 79906
rect 173222 79898 173250 80036
rect 173210 79892 173262 79898
rect 173210 79834 173262 79840
rect 172946 79784 173020 79812
rect 172854 79716 172928 79744
rect 172762 79614 172836 79642
rect 172704 79484 172756 79490
rect 172704 79426 172756 79432
rect 172716 78985 172744 79426
rect 172702 78976 172758 78985
rect 172702 78911 172758 78920
rect 172808 76838 172836 79614
rect 172900 79014 172928 79716
rect 172888 79008 172940 79014
rect 172888 78950 172940 78956
rect 172992 78198 173020 79784
rect 173070 79792 173126 79801
rect 173314 79744 173342 80036
rect 173406 79830 173434 80036
rect 173394 79824 173446 79830
rect 173394 79766 173446 79772
rect 173498 79778 173526 80036
rect 173590 79898 173618 80036
rect 173578 79892 173630 79898
rect 173578 79834 173630 79840
rect 173498 79750 173572 79778
rect 173070 79727 173126 79736
rect 173084 78606 173112 79727
rect 173176 79716 173342 79744
rect 173072 78600 173124 78606
rect 173072 78542 173124 78548
rect 172980 78192 173032 78198
rect 172980 78134 173032 78140
rect 173070 78160 173126 78169
rect 173070 78095 173126 78104
rect 172796 76832 172848 76838
rect 172796 76774 172848 76780
rect 173084 71233 173112 78095
rect 173176 75585 173204 79716
rect 173440 79688 173492 79694
rect 173440 79630 173492 79636
rect 173256 79620 173308 79626
rect 173256 79562 173308 79568
rect 173162 75576 173218 75585
rect 173162 75511 173218 75520
rect 173070 71224 173126 71233
rect 173070 71159 173126 71168
rect 172612 70372 172664 70378
rect 172612 70314 172664 70320
rect 172060 70100 172112 70106
rect 172060 70042 172112 70048
rect 171968 69896 172020 69902
rect 171968 69838 172020 69844
rect 171876 68876 171928 68882
rect 171876 68818 171928 68824
rect 171888 67998 171916 68818
rect 171968 68536 172020 68542
rect 171968 68478 172020 68484
rect 171980 68066 172008 68478
rect 172060 68400 172112 68406
rect 172058 68368 172060 68377
rect 172112 68368 172114 68377
rect 172058 68303 172114 68312
rect 171968 68060 172020 68066
rect 171968 68002 172020 68008
rect 171876 67992 171928 67998
rect 171876 67934 171928 67940
rect 171876 64864 171928 64870
rect 171876 64806 171928 64812
rect 171888 64598 171916 64806
rect 171876 64592 171928 64598
rect 171876 64534 171928 64540
rect 171888 26314 171916 64534
rect 173268 64530 173296 79562
rect 173348 75948 173400 75954
rect 173348 75890 173400 75896
rect 173360 69834 173388 75890
rect 173452 71262 173480 79630
rect 173544 79626 173572 79750
rect 173682 79744 173710 80036
rect 173774 79966 173802 80036
rect 173762 79960 173814 79966
rect 173762 79902 173814 79908
rect 173866 79812 173894 80036
rect 173958 79971 173986 80036
rect 173944 79962 174000 79971
rect 173944 79897 174000 79906
rect 174050 79898 174078 80036
rect 174142 79898 174170 80036
rect 174038 79892 174090 79898
rect 174038 79834 174090 79840
rect 174130 79892 174182 79898
rect 174130 79834 174182 79840
rect 173820 79784 173894 79812
rect 173682 79716 173756 79744
rect 173532 79620 173584 79626
rect 173532 79562 173584 79568
rect 173624 79620 173676 79626
rect 173624 79562 173676 79568
rect 173532 79484 173584 79490
rect 173532 79426 173584 79432
rect 173544 79354 173572 79426
rect 173532 79348 173584 79354
rect 173532 79290 173584 79296
rect 173532 77920 173584 77926
rect 173532 77862 173584 77868
rect 173440 71256 173492 71262
rect 173440 71198 173492 71204
rect 173348 69828 173400 69834
rect 173348 69770 173400 69776
rect 173544 68377 173572 77862
rect 173636 77042 173664 79562
rect 173624 77036 173676 77042
rect 173624 76978 173676 76984
rect 173728 75954 173756 79716
rect 173716 75948 173768 75954
rect 173716 75890 173768 75896
rect 173820 75721 173848 79784
rect 174234 79744 174262 80036
rect 174188 79716 174262 79744
rect 173900 79688 173952 79694
rect 173900 79630 173952 79636
rect 173806 75712 173862 75721
rect 173806 75647 173862 75656
rect 173912 73001 173940 79630
rect 173992 79620 174044 79626
rect 173992 79562 174044 79568
rect 173898 72992 173954 73001
rect 173898 72927 173954 72936
rect 173808 71732 173860 71738
rect 173808 71674 173860 71680
rect 173820 70446 173848 71674
rect 173808 70440 173860 70446
rect 173808 70382 173860 70388
rect 173530 68368 173586 68377
rect 173530 68303 173586 68312
rect 173820 65890 173848 70382
rect 173900 69692 173952 69698
rect 173900 69634 173952 69640
rect 173808 65884 173860 65890
rect 173808 65826 173860 65832
rect 173256 64524 173308 64530
rect 173256 64466 173308 64472
rect 173808 64524 173860 64530
rect 173808 64466 173860 64472
rect 171876 26308 171928 26314
rect 171876 26250 171928 26256
rect 173820 25634 173848 64466
rect 173808 25628 173860 25634
rect 173808 25570 173860 25576
rect 173912 16574 173940 69634
rect 174004 64666 174032 79562
rect 174084 79008 174136 79014
rect 174084 78950 174136 78956
rect 174096 78674 174124 78950
rect 174084 78668 174136 78674
rect 174084 78610 174136 78616
rect 174084 75268 174136 75274
rect 174084 75210 174136 75216
rect 174096 67386 174124 75210
rect 174188 70038 174216 79716
rect 174326 79472 174354 80036
rect 174418 79540 174446 80036
rect 174510 79830 174538 80036
rect 174602 79830 174630 80036
rect 174498 79824 174550 79830
rect 174498 79766 174550 79772
rect 174590 79824 174642 79830
rect 174590 79766 174642 79772
rect 174694 79744 174722 80036
rect 174786 79812 174814 80036
rect 174878 79966 174906 80036
rect 174970 79966 174998 80036
rect 174866 79960 174918 79966
rect 174866 79902 174918 79908
rect 174958 79960 175010 79966
rect 174958 79902 175010 79908
rect 174912 79824 174964 79830
rect 174786 79801 174860 79812
rect 174786 79792 174874 79801
rect 174786 79784 174818 79792
rect 174694 79716 174768 79744
rect 174912 79766 174964 79772
rect 175062 79778 175090 80036
rect 175154 79898 175182 80036
rect 175142 79892 175194 79898
rect 175142 79834 175194 79840
rect 175246 79778 175274 80036
rect 175338 79898 175366 80036
rect 175430 79966 175458 80036
rect 175418 79960 175470 79966
rect 175418 79902 175470 79908
rect 175326 79892 175378 79898
rect 175326 79834 175378 79840
rect 175522 79830 175550 80036
rect 175614 79830 175642 80036
rect 174818 79727 174874 79736
rect 174544 79620 174596 79626
rect 174544 79562 174596 79568
rect 174418 79512 174492 79540
rect 174326 79444 174400 79472
rect 174372 75274 174400 79444
rect 174464 75914 174492 79512
rect 174556 78010 174584 79562
rect 174740 79393 174768 79716
rect 174820 79688 174872 79694
rect 174820 79630 174872 79636
rect 174726 79384 174782 79393
rect 174726 79319 174782 79328
rect 174832 78282 174860 79630
rect 174924 79218 174952 79766
rect 175062 79750 175136 79778
rect 175004 79688 175056 79694
rect 175004 79630 175056 79636
rect 174912 79212 174964 79218
rect 174912 79154 174964 79160
rect 174832 78254 174952 78282
rect 174728 78192 174780 78198
rect 174726 78160 174728 78169
rect 174820 78192 174872 78198
rect 174780 78160 174782 78169
rect 174820 78134 174872 78140
rect 174726 78095 174782 78104
rect 174556 77982 174768 78010
rect 174634 76528 174690 76537
rect 174634 76463 174690 76472
rect 174464 75886 174584 75914
rect 174556 75478 174584 75886
rect 174544 75472 174596 75478
rect 174544 75414 174596 75420
rect 174360 75268 174412 75274
rect 174360 75210 174412 75216
rect 174544 75132 174596 75138
rect 174544 75074 174596 75080
rect 174176 70032 174228 70038
rect 174176 69974 174228 69980
rect 174084 67380 174136 67386
rect 174084 67322 174136 67328
rect 173992 64660 174044 64666
rect 173992 64602 174044 64608
rect 173912 16546 174492 16574
rect 171784 4888 171836 4894
rect 171784 4830 171836 4836
rect 174464 490 174492 16546
rect 174556 3670 174584 75074
rect 174648 67425 174676 76463
rect 174740 71398 174768 77982
rect 174728 71392 174780 71398
rect 174728 71334 174780 71340
rect 174634 67416 174690 67425
rect 174634 67351 174690 67360
rect 174832 61402 174860 78134
rect 174924 71738 174952 78254
rect 175016 78198 175044 79630
rect 175108 78441 175136 79750
rect 175200 79750 175274 79778
rect 175510 79824 175562 79830
rect 175510 79766 175562 79772
rect 175602 79824 175654 79830
rect 175602 79766 175654 79772
rect 175706 79778 175734 80036
rect 175798 79898 175826 80036
rect 175890 79966 175918 80036
rect 175982 79971 176010 80036
rect 175878 79960 175930 79966
rect 175878 79902 175930 79908
rect 175968 79962 176024 79971
rect 175786 79892 175838 79898
rect 175968 79897 176024 79906
rect 175786 79834 175838 79840
rect 176074 79778 176102 80036
rect 176166 79966 176194 80036
rect 176258 79966 176286 80036
rect 176350 79971 176378 80036
rect 176154 79960 176206 79966
rect 176154 79902 176206 79908
rect 176246 79960 176298 79966
rect 176246 79902 176298 79908
rect 176336 79962 176392 79971
rect 176442 79966 176470 80036
rect 176336 79897 176392 79906
rect 176430 79960 176482 79966
rect 176430 79902 176482 79908
rect 176200 79824 176252 79830
rect 175372 79756 175424 79762
rect 175094 78432 175150 78441
rect 175094 78367 175150 78376
rect 175004 78192 175056 78198
rect 175004 78134 175056 78140
rect 175200 76158 175228 79750
rect 175706 79750 175780 79778
rect 175372 79698 175424 79704
rect 175280 79688 175332 79694
rect 175280 79630 175332 79636
rect 175188 76152 175240 76158
rect 175188 76094 175240 76100
rect 175292 71738 175320 79630
rect 175384 79393 175412 79698
rect 175464 79688 175516 79694
rect 175464 79630 175516 79636
rect 175648 79688 175700 79694
rect 175648 79630 175700 79636
rect 175370 79384 175426 79393
rect 175370 79319 175426 79328
rect 175372 79280 175424 79286
rect 175372 79222 175424 79228
rect 175384 76974 175412 79222
rect 175372 76968 175424 76974
rect 175372 76910 175424 76916
rect 174912 71732 174964 71738
rect 174912 71674 174964 71680
rect 175280 71732 175332 71738
rect 175280 71674 175332 71680
rect 175476 64870 175504 79630
rect 175556 79280 175608 79286
rect 175556 79222 175608 79228
rect 175568 75750 175596 79222
rect 175556 75744 175608 75750
rect 175556 75686 175608 75692
rect 175660 72622 175688 79630
rect 175752 74458 175780 79750
rect 175832 79756 175884 79762
rect 176074 79750 176148 79778
rect 176534 79812 176562 80036
rect 176200 79766 176252 79772
rect 176488 79784 176562 79812
rect 175832 79698 175884 79704
rect 175844 75682 175872 79698
rect 176016 79688 176068 79694
rect 176016 79630 176068 79636
rect 175924 79552 175976 79558
rect 175924 79494 175976 79500
rect 175936 78538 175964 79494
rect 175924 78532 175976 78538
rect 175924 78474 175976 78480
rect 176028 75857 176056 79630
rect 176120 77246 176148 79750
rect 176108 77240 176160 77246
rect 176108 77182 176160 77188
rect 176014 75848 176070 75857
rect 176014 75783 176070 75792
rect 175832 75676 175884 75682
rect 175832 75618 175884 75624
rect 175844 74534 175872 75618
rect 176212 75313 176240 79766
rect 176292 79620 176344 79626
rect 176292 79562 176344 79568
rect 176304 79286 176332 79562
rect 176488 79286 176516 79784
rect 176626 79744 176654 80036
rect 176718 79898 176746 80036
rect 176810 79898 176838 80036
rect 176706 79892 176758 79898
rect 176706 79834 176758 79840
rect 176798 79892 176850 79898
rect 176798 79834 176850 79840
rect 176580 79716 176654 79744
rect 176750 79792 176806 79801
rect 176750 79727 176806 79736
rect 176902 79744 176930 80036
rect 176994 79898 177022 80036
rect 177086 79898 177114 80036
rect 177178 79898 177206 80036
rect 176982 79892 177034 79898
rect 176982 79834 177034 79840
rect 177074 79892 177126 79898
rect 177074 79834 177126 79840
rect 177166 79892 177218 79898
rect 177166 79834 177218 79840
rect 177270 79801 177298 80036
rect 177256 79792 177312 79801
rect 176292 79280 176344 79286
rect 176292 79222 176344 79228
rect 176476 79280 176528 79286
rect 176476 79222 176528 79228
rect 176476 76628 176528 76634
rect 176476 76570 176528 76576
rect 176198 75304 176254 75313
rect 176198 75239 176254 75248
rect 175844 74506 176056 74534
rect 175740 74452 175792 74458
rect 175740 74394 175792 74400
rect 175648 72616 175700 72622
rect 175648 72558 175700 72564
rect 175464 64864 175516 64870
rect 175464 64806 175516 64812
rect 175924 64864 175976 64870
rect 175924 64806 175976 64812
rect 175188 64660 175240 64666
rect 175188 64602 175240 64608
rect 174820 61396 174872 61402
rect 174820 61338 174872 61344
rect 175200 26926 175228 64602
rect 175188 26920 175240 26926
rect 175188 26862 175240 26868
rect 175936 9110 175964 64806
rect 176028 10402 176056 74506
rect 176108 71732 176160 71738
rect 176108 71674 176160 71680
rect 176120 71058 176148 71674
rect 176108 71052 176160 71058
rect 176108 70994 176160 71000
rect 176120 55962 176148 70994
rect 176488 68241 176516 76570
rect 176580 71670 176608 79716
rect 176660 79620 176712 79626
rect 176660 79562 176712 79568
rect 176568 71664 176620 71670
rect 176568 71606 176620 71612
rect 176474 68232 176530 68241
rect 176474 68167 176530 68176
rect 176672 67522 176700 79562
rect 176764 79014 176792 79727
rect 176902 79716 176976 79744
rect 177256 79727 177312 79736
rect 176948 79642 176976 79716
rect 177362 79676 177390 80036
rect 177454 79744 177482 80036
rect 177546 79914 177574 80036
rect 177638 80016 177666 80036
rect 177638 79988 177712 80016
rect 177546 79886 177620 79914
rect 177454 79716 177528 79744
rect 177316 79648 177390 79676
rect 176948 79626 177160 79642
rect 176948 79620 177172 79626
rect 176948 79614 177120 79620
rect 177120 79562 177172 79568
rect 176844 79552 176896 79558
rect 176844 79494 176896 79500
rect 177028 79552 177080 79558
rect 177028 79494 177080 79500
rect 176752 79008 176804 79014
rect 176752 78950 176804 78956
rect 176752 75948 176804 75954
rect 176752 75890 176804 75896
rect 176764 70242 176792 75890
rect 176752 70236 176804 70242
rect 176752 70178 176804 70184
rect 176856 69698 176884 79494
rect 177040 70990 177068 79494
rect 177316 76809 177344 79648
rect 177396 79552 177448 79558
rect 177396 79494 177448 79500
rect 177408 78266 177436 79494
rect 177396 78260 177448 78266
rect 177396 78202 177448 78208
rect 177302 76800 177358 76809
rect 177500 76770 177528 79716
rect 177592 78577 177620 79886
rect 177578 78568 177634 78577
rect 177578 78503 177634 78512
rect 177302 76735 177358 76744
rect 177488 76764 177540 76770
rect 177488 76706 177540 76712
rect 177684 75954 177712 79988
rect 177776 79898 177804 80174
rect 177868 79966 177896 80650
rect 177960 80617 177988 80650
rect 177946 80608 178002 80617
rect 177946 80543 178002 80552
rect 179604 80504 179656 80510
rect 179234 80472 179290 80481
rect 178132 80436 178184 80442
rect 179604 80446 179656 80452
rect 179234 80407 179290 80416
rect 178132 80378 178184 80384
rect 178040 80300 178092 80306
rect 178040 80242 178092 80248
rect 177856 79960 177908 79966
rect 177856 79902 177908 79908
rect 177946 79928 178002 79937
rect 177764 79892 177816 79898
rect 177946 79863 178002 79872
rect 177764 79834 177816 79840
rect 177960 76537 177988 79863
rect 178052 79762 178080 80242
rect 178040 79756 178092 79762
rect 178040 79698 178092 79704
rect 178144 78946 178172 80378
rect 178960 80232 179012 80238
rect 178960 80174 179012 80180
rect 178132 78940 178184 78946
rect 178132 78882 178184 78888
rect 177946 76528 178002 76537
rect 177946 76463 178002 76472
rect 177948 76152 178000 76158
rect 177948 76094 178000 76100
rect 177672 75948 177724 75954
rect 177672 75890 177724 75896
rect 177960 75138 177988 76094
rect 178972 75449 179000 80174
rect 179248 80102 179276 80407
rect 179236 80096 179288 80102
rect 179616 80073 179644 80446
rect 179236 80038 179288 80044
rect 179602 80064 179658 80073
rect 182836 80034 182864 80650
rect 188344 80640 188396 80646
rect 186318 80608 186374 80617
rect 188344 80582 188396 80588
rect 186318 80543 186374 80552
rect 186964 80572 187016 80578
rect 185582 80472 185638 80481
rect 185582 80407 185638 80416
rect 179602 79999 179658 80008
rect 182824 80028 182876 80034
rect 182824 79970 182876 79976
rect 183928 80028 183980 80034
rect 183928 79970 183980 79976
rect 179052 79892 179104 79898
rect 179052 79834 179104 79840
rect 179064 77761 179092 79834
rect 179788 79620 179840 79626
rect 179788 79562 179840 79568
rect 179050 77752 179106 77761
rect 179050 77687 179106 77696
rect 179800 76634 179828 79562
rect 181352 79144 181404 79150
rect 181352 79086 181404 79092
rect 181364 78742 181392 79086
rect 181444 79076 181496 79082
rect 181444 79018 181496 79024
rect 181456 78962 181484 79018
rect 181628 79008 181680 79014
rect 181456 78956 181628 78962
rect 181456 78950 181680 78956
rect 181456 78934 181668 78950
rect 181352 78736 181404 78742
rect 181352 78678 181404 78684
rect 182180 78736 182232 78742
rect 182180 78678 182232 78684
rect 181812 78260 181864 78266
rect 181812 78202 181864 78208
rect 180524 78056 180576 78062
rect 180524 77998 180576 78004
rect 180708 78056 180760 78062
rect 180708 77998 180760 78004
rect 180340 77988 180392 77994
rect 180340 77930 180392 77936
rect 179970 77888 180026 77897
rect 179970 77823 180026 77832
rect 179788 76628 179840 76634
rect 179788 76570 179840 76576
rect 178958 75440 179014 75449
rect 178958 75375 179014 75384
rect 177948 75132 178000 75138
rect 177948 75074 178000 75080
rect 179984 74934 180012 77823
rect 180352 76362 180380 77930
rect 180340 76356 180392 76362
rect 180340 76298 180392 76304
rect 180536 75342 180564 77998
rect 180720 76294 180748 77998
rect 180708 76288 180760 76294
rect 180708 76230 180760 76236
rect 180524 75336 180576 75342
rect 180524 75278 180576 75284
rect 179972 74928 180024 74934
rect 179972 74870 180024 74876
rect 177028 70984 177080 70990
rect 177028 70926 177080 70932
rect 177040 70394 177068 70926
rect 180536 70394 180564 75278
rect 181444 75200 181496 75206
rect 181444 75142 181496 75148
rect 181456 74361 181484 75142
rect 181824 74866 181852 78202
rect 182192 78169 182220 78678
rect 183940 78441 183968 79970
rect 185596 79966 185624 80407
rect 185584 79960 185636 79966
rect 185584 79902 185636 79908
rect 186332 79121 186360 80543
rect 186964 80514 187016 80520
rect 186318 79112 186374 79121
rect 186318 79047 186374 79056
rect 183926 78432 183982 78441
rect 183926 78367 183982 78376
rect 184202 78432 184258 78441
rect 184202 78367 184258 78376
rect 186318 78432 186374 78441
rect 186318 78367 186374 78376
rect 182178 78160 182234 78169
rect 182088 78124 182140 78130
rect 182178 78095 182234 78104
rect 182916 78124 182968 78130
rect 182088 78066 182140 78072
rect 182916 78066 182968 78072
rect 181812 74860 181864 74866
rect 181812 74802 181864 74808
rect 181442 74352 181498 74361
rect 181442 74287 181498 74296
rect 182100 73642 182128 78066
rect 182824 77920 182876 77926
rect 182824 77862 182876 77868
rect 182180 73908 182232 73914
rect 182180 73850 182232 73856
rect 182088 73636 182140 73642
rect 182088 73578 182140 73584
rect 177040 70366 177344 70394
rect 180536 70366 180748 70394
rect 176844 69692 176896 69698
rect 176844 69634 176896 69640
rect 176660 67516 176712 67522
rect 176660 67458 176712 67464
rect 176108 55956 176160 55962
rect 176108 55898 176160 55904
rect 177316 33046 177344 70366
rect 177304 33040 177356 33046
rect 177304 32982 177356 32988
rect 180720 20670 180748 70366
rect 180708 20664 180760 20670
rect 180708 20606 180760 20612
rect 182100 12442 182128 73578
rect 182192 73166 182220 73850
rect 182180 73160 182232 73166
rect 182180 73102 182232 73108
rect 182836 68950 182864 77862
rect 182824 68944 182876 68950
rect 182824 68886 182876 68892
rect 182928 68202 182956 78066
rect 183468 73160 183520 73166
rect 183468 73102 183520 73108
rect 182916 68196 182968 68202
rect 182916 68138 182968 68144
rect 182180 62892 182232 62898
rect 182180 62834 182232 62840
rect 182192 16574 182220 62834
rect 183480 49706 183508 73102
rect 183468 49700 183520 49706
rect 183468 49642 183520 49648
rect 184216 24818 184244 78367
rect 185584 72480 185636 72486
rect 185584 72422 185636 72428
rect 185596 41410 185624 72422
rect 186332 62014 186360 78367
rect 186976 70281 187004 80514
rect 187056 80504 187108 80510
rect 187056 80446 187108 80452
rect 187068 70922 187096 80446
rect 187056 70916 187108 70922
rect 187056 70858 187108 70864
rect 186962 70272 187018 70281
rect 186962 70207 187018 70216
rect 188356 65822 188384 80582
rect 188434 80472 188490 80481
rect 188434 80407 188490 80416
rect 188448 74497 188476 80407
rect 188632 80209 188660 80990
rect 188618 80200 188674 80209
rect 188618 80135 188674 80144
rect 188724 78334 188752 193190
rect 188804 191616 188856 191622
rect 188804 191558 188856 191564
rect 188816 78674 188844 191558
rect 188896 184000 188948 184006
rect 188896 183942 188948 183948
rect 188908 145042 188936 183942
rect 188896 145036 188948 145042
rect 188896 144978 188948 144984
rect 189000 144922 189028 199718
rect 189264 198348 189316 198354
rect 189264 198290 189316 198296
rect 189172 198280 189224 198286
rect 189172 198222 189224 198228
rect 189078 195256 189134 195265
rect 189078 195191 189134 195200
rect 189092 194857 189120 195191
rect 189078 194848 189134 194857
rect 189078 194783 189134 194792
rect 189080 189644 189132 189650
rect 189080 189586 189132 189592
rect 188908 144894 189028 144922
rect 188908 140049 188936 144894
rect 188988 142452 189040 142458
rect 188988 142394 189040 142400
rect 188894 140040 188950 140049
rect 188894 139975 188950 139984
rect 188896 139868 188948 139874
rect 188896 139810 188948 139816
rect 188908 138014 188936 139810
rect 189000 138718 189028 142394
rect 188988 138712 189040 138718
rect 188988 138654 189040 138660
rect 188908 137986 189028 138014
rect 189000 137834 189028 137986
rect 188988 137828 189040 137834
rect 188988 137770 189040 137776
rect 188986 91216 189042 91225
rect 188986 91151 189042 91160
rect 188896 81728 188948 81734
rect 188896 81670 188948 81676
rect 188804 78668 188856 78674
rect 188804 78610 188856 78616
rect 188908 78402 188936 81670
rect 188896 78396 188948 78402
rect 188896 78338 188948 78344
rect 188712 78328 188764 78334
rect 188712 78270 188764 78276
rect 188434 74488 188490 74497
rect 188434 74423 188490 74432
rect 189000 66201 189028 91151
rect 188986 66192 189042 66201
rect 188986 66127 189042 66136
rect 188344 65816 188396 65822
rect 188344 65758 188396 65764
rect 189092 64190 189120 189586
rect 189184 84862 189212 198222
rect 189276 186046 189304 198290
rect 189460 192846 189488 700062
rect 189632 265804 189684 265810
rect 189632 265746 189684 265752
rect 189540 264988 189592 264994
rect 189540 264930 189592 264936
rect 189448 192840 189500 192846
rect 189448 192782 189500 192788
rect 189356 189576 189408 189582
rect 189356 189518 189408 189524
rect 189264 186040 189316 186046
rect 189264 185982 189316 185988
rect 189264 181824 189316 181830
rect 189264 181766 189316 181772
rect 189172 84856 189224 84862
rect 189172 84798 189224 84804
rect 189172 82136 189224 82142
rect 189172 82078 189224 82084
rect 189184 79490 189212 82078
rect 189172 79484 189224 79490
rect 189172 79426 189224 79432
rect 189080 64184 189132 64190
rect 189080 64126 189132 64132
rect 189092 63986 189120 64126
rect 189276 64054 189304 181766
rect 189368 72690 189396 189518
rect 189448 182096 189500 182102
rect 189448 182038 189500 182044
rect 189356 72684 189408 72690
rect 189356 72626 189408 72632
rect 189460 65686 189488 182038
rect 189552 144702 189580 264930
rect 189644 197266 189672 265746
rect 189736 199617 189764 700266
rect 191748 419552 191800 419558
rect 191748 419494 191800 419500
rect 189816 386436 189868 386442
rect 189816 386378 189868 386384
rect 189722 199608 189778 199617
rect 189828 199578 189856 386378
rect 189908 367124 189960 367130
rect 189908 367066 189960 367072
rect 189722 199543 189778 199552
rect 189816 199572 189868 199578
rect 189816 199514 189868 199520
rect 189920 198762 189948 367066
rect 191656 272536 191708 272542
rect 191656 272478 191708 272484
rect 191668 271930 191696 272478
rect 190460 271924 190512 271930
rect 190460 271866 190512 271872
rect 191656 271924 191708 271930
rect 191656 271866 191708 271872
rect 190000 265940 190052 265946
rect 190000 265882 190052 265888
rect 189908 198756 189960 198762
rect 189908 198698 189960 198704
rect 190012 197577 190040 265882
rect 190092 225004 190144 225010
rect 190092 224946 190144 224952
rect 190104 199034 190132 224946
rect 190092 199028 190144 199034
rect 190092 198970 190144 198976
rect 189998 197568 190054 197577
rect 190054 197526 190132 197554
rect 189998 197503 190054 197512
rect 189632 197260 189684 197266
rect 189632 197202 189684 197208
rect 189906 195256 189962 195265
rect 189906 195191 189962 195200
rect 189632 194268 189684 194274
rect 189632 194210 189684 194216
rect 189540 144696 189592 144702
rect 189540 144638 189592 144644
rect 189540 140072 189592 140078
rect 189540 140014 189592 140020
rect 189448 65680 189500 65686
rect 189448 65622 189500 65628
rect 189264 64048 189316 64054
rect 189264 63990 189316 63996
rect 189080 63980 189132 63986
rect 189080 63922 189132 63928
rect 186320 62008 186372 62014
rect 186320 61950 186372 61956
rect 189552 57866 189580 140014
rect 189644 85082 189672 194210
rect 189724 192432 189776 192438
rect 189724 192374 189776 192380
rect 189736 85202 189764 192374
rect 189816 147348 189868 147354
rect 189816 147290 189868 147296
rect 189828 89714 189856 147290
rect 189920 136649 189948 195191
rect 190000 194540 190052 194546
rect 190000 194482 190052 194488
rect 190012 194274 190040 194482
rect 190000 194268 190052 194274
rect 190000 194210 190052 194216
rect 190104 194206 190132 197526
rect 190092 194200 190144 194206
rect 190092 194142 190144 194148
rect 190472 142361 190500 271866
rect 190828 263152 190880 263158
rect 190828 263094 190880 263100
rect 190644 262812 190696 262818
rect 190644 262754 190696 262760
rect 190552 260228 190604 260234
rect 190552 260170 190604 260176
rect 190564 204950 190592 260170
rect 190552 204944 190604 204950
rect 190552 204886 190604 204892
rect 190552 200252 190604 200258
rect 190552 200194 190604 200200
rect 190564 199170 190592 200194
rect 190552 199164 190604 199170
rect 190552 199106 190604 199112
rect 190552 184136 190604 184142
rect 190552 184078 190604 184084
rect 190458 142352 190514 142361
rect 190458 142287 190514 142296
rect 190460 140004 190512 140010
rect 190460 139946 190512 139952
rect 189906 136640 189962 136649
rect 189906 136575 189962 136584
rect 189828 89686 189948 89714
rect 189724 85196 189776 85202
rect 189724 85138 189776 85144
rect 189644 85054 189856 85082
rect 189724 84924 189776 84930
rect 189724 84866 189776 84872
rect 189632 84856 189684 84862
rect 189632 84798 189684 84804
rect 189644 77217 189672 84798
rect 189736 78198 189764 84866
rect 189828 80054 189856 85054
rect 189920 80646 189948 89686
rect 189998 81424 190054 81433
rect 189998 81359 190054 81368
rect 189908 80640 189960 80646
rect 189908 80582 189960 80588
rect 190012 80481 190040 81359
rect 189998 80472 190054 80481
rect 189998 80407 190054 80416
rect 189828 80026 189948 80054
rect 189724 78192 189776 78198
rect 189724 78134 189776 78140
rect 189920 77722 189948 80026
rect 189908 77716 189960 77722
rect 189908 77658 189960 77664
rect 189630 77208 189686 77217
rect 189630 77143 189686 77152
rect 190472 72758 190500 139946
rect 190460 72752 190512 72758
rect 190460 72694 190512 72700
rect 190460 68264 190512 68270
rect 190460 68206 190512 68212
rect 189080 57860 189132 57866
rect 189080 57802 189132 57808
rect 189540 57860 189592 57866
rect 189540 57802 189592 57808
rect 189092 57254 189120 57802
rect 189080 57248 189132 57254
rect 189080 57190 189132 57196
rect 185584 41404 185636 41410
rect 185584 41346 185636 41352
rect 184204 24812 184256 24818
rect 184204 24754 184256 24760
rect 182192 16546 182496 16574
rect 182088 12436 182140 12442
rect 182088 12378 182140 12384
rect 176016 10396 176068 10402
rect 176016 10338 176068 10344
rect 175924 9104 175976 9110
rect 175924 9046 175976 9052
rect 174544 3664 174596 3670
rect 174544 3606 174596 3612
rect 179052 3596 179104 3602
rect 179052 3538 179104 3544
rect 171294 354 171406 480
rect 174464 462 174860 490
rect 179064 480 179092 3538
rect 171152 326 171406 354
rect 174832 354 174860 462
rect 175158 354 175270 480
rect 174832 326 175270 354
rect 171294 -960 171406 326
rect 175158 -960 175270 326
rect 179022 -960 179134 480
rect 182468 354 182496 16546
rect 186780 3664 186832 3670
rect 186780 3606 186832 3612
rect 186792 480 186820 3606
rect 182886 354 182998 480
rect 182468 326 182998 354
rect 182886 -960 182998 326
rect 186750 -960 186862 480
rect 190472 354 190500 68206
rect 190564 61946 190592 184078
rect 190656 141846 190684 262754
rect 190736 262404 190788 262410
rect 190736 262346 190788 262352
rect 190748 141914 190776 262346
rect 190840 144634 190868 263094
rect 191104 262744 191156 262750
rect 191104 262686 191156 262692
rect 190920 204944 190972 204950
rect 190920 204886 190972 204892
rect 190932 194478 190960 204886
rect 190920 194472 190972 194478
rect 190920 194414 190972 194420
rect 191012 190324 191064 190330
rect 191012 190266 191064 190272
rect 190920 190120 190972 190126
rect 190920 190062 190972 190068
rect 190828 144628 190880 144634
rect 190828 144570 190880 144576
rect 190736 141908 190788 141914
rect 190736 141850 190788 141856
rect 190644 141840 190696 141846
rect 190644 141782 190696 141788
rect 190656 141506 190684 141782
rect 190644 141500 190696 141506
rect 190644 141442 190696 141448
rect 190828 141432 190880 141438
rect 190828 141374 190880 141380
rect 190644 141364 190696 141370
rect 190644 141306 190696 141312
rect 190552 61940 190604 61946
rect 190552 61882 190604 61888
rect 190656 48278 190684 141306
rect 190736 140684 190788 140690
rect 190736 140626 190788 140632
rect 190748 73710 190776 140626
rect 190840 80034 190868 141374
rect 190828 80028 190880 80034
rect 190828 79970 190880 79976
rect 190736 73704 190788 73710
rect 190736 73646 190788 73652
rect 190932 72962 190960 190062
rect 191024 74526 191052 190266
rect 191116 143682 191144 262686
rect 191656 253972 191708 253978
rect 191656 253914 191708 253920
rect 191196 241528 191248 241534
rect 191196 241470 191248 241476
rect 191208 200705 191236 241470
rect 191668 204218 191696 253914
rect 191484 204190 191696 204218
rect 191484 201550 191512 204190
rect 191760 203402 191788 419494
rect 191668 203374 191788 203402
rect 191472 201544 191524 201550
rect 191472 201486 191524 201492
rect 191194 200696 191250 200705
rect 191194 200631 191250 200640
rect 191668 200258 191696 203374
rect 191748 201544 191800 201550
rect 191748 201486 191800 201492
rect 191760 200666 191788 201486
rect 191748 200660 191800 200666
rect 191748 200602 191800 200608
rect 191656 200252 191708 200258
rect 191656 200194 191708 200200
rect 191196 196036 191248 196042
rect 191196 195978 191248 195984
rect 191208 177886 191236 195978
rect 191852 194546 191880 700402
rect 193220 700392 193272 700398
rect 193220 700334 193272 700340
rect 192484 535492 192536 535498
rect 192484 535434 192536 535440
rect 192392 260908 192444 260914
rect 192392 260850 192444 260856
rect 192300 260160 192352 260166
rect 192300 260102 192352 260108
rect 192024 260092 192076 260098
rect 192024 260034 192076 260040
rect 191932 197124 191984 197130
rect 191932 197066 191984 197072
rect 191840 194540 191892 194546
rect 191840 194482 191892 194488
rect 191944 182238 191972 197066
rect 191932 182232 191984 182238
rect 191932 182174 191984 182180
rect 191196 177880 191248 177886
rect 191196 177822 191248 177828
rect 191932 160744 191984 160750
rect 191932 160686 191984 160692
rect 191840 144288 191892 144294
rect 191840 144230 191892 144236
rect 191104 143676 191156 143682
rect 191104 143618 191156 143624
rect 191116 142866 191144 143618
rect 191104 142860 191156 142866
rect 191104 142802 191156 142808
rect 191196 141704 191248 141710
rect 191196 141646 191248 141652
rect 191104 141636 191156 141642
rect 191104 141578 191156 141584
rect 191116 80510 191144 141578
rect 191208 82793 191236 141646
rect 191288 91112 191340 91118
rect 191288 91054 191340 91060
rect 191194 82784 191250 82793
rect 191194 82719 191250 82728
rect 191104 80504 191156 80510
rect 191104 80446 191156 80452
rect 191012 74520 191064 74526
rect 191012 74462 191064 74468
rect 190920 72956 190972 72962
rect 190920 72898 190972 72904
rect 191300 64122 191328 91054
rect 191748 72956 191800 72962
rect 191748 72898 191800 72904
rect 191760 72486 191788 72898
rect 191748 72480 191800 72486
rect 191748 72422 191800 72428
rect 191852 68746 191880 144230
rect 191944 75886 191972 160686
rect 192036 143342 192064 260034
rect 192208 259820 192260 259826
rect 192208 259762 192260 259768
rect 192116 259548 192168 259554
rect 192116 259490 192168 259496
rect 192024 143336 192076 143342
rect 192024 143278 192076 143284
rect 192128 143041 192156 259490
rect 192114 143032 192170 143041
rect 192114 142967 192170 142976
rect 192128 142866 192156 142967
rect 192220 142934 192248 259762
rect 192312 197334 192340 260102
rect 192300 197328 192352 197334
rect 192300 197270 192352 197276
rect 192300 189848 192352 189854
rect 192300 189790 192352 189796
rect 192208 142928 192260 142934
rect 192208 142870 192260 142876
rect 192116 142860 192168 142866
rect 192116 142802 192168 142808
rect 192116 142044 192168 142050
rect 192116 141986 192168 141992
rect 191932 75880 191984 75886
rect 191932 75822 191984 75828
rect 191840 68740 191892 68746
rect 191840 68682 191892 68688
rect 192128 65958 192156 141986
rect 192206 139360 192262 139369
rect 192206 139295 192262 139304
rect 192220 67017 192248 139295
rect 192312 74322 192340 189790
rect 192404 145518 192432 260850
rect 192496 199782 192524 535434
rect 192576 503736 192628 503742
rect 192576 503678 192628 503684
rect 192588 264450 192616 503678
rect 192576 264444 192628 264450
rect 192576 264386 192628 264392
rect 192852 262540 192904 262546
rect 192852 262482 192904 262488
rect 192576 260976 192628 260982
rect 192576 260918 192628 260924
rect 192588 251190 192616 260918
rect 192576 251184 192628 251190
rect 192576 251126 192628 251132
rect 192484 199776 192536 199782
rect 192484 199718 192536 199724
rect 192576 197192 192628 197198
rect 192576 197134 192628 197140
rect 192484 189984 192536 189990
rect 192484 189926 192536 189932
rect 192392 145512 192444 145518
rect 192392 145454 192444 145460
rect 192390 143576 192446 143585
rect 192390 143511 192446 143520
rect 192404 142934 192432 143511
rect 192392 142928 192444 142934
rect 192392 142870 192444 142876
rect 192392 140752 192444 140758
rect 192392 140694 192444 140700
rect 192300 74316 192352 74322
rect 192300 74258 192352 74264
rect 192404 72418 192432 140694
rect 192496 76906 192524 189926
rect 192588 162178 192616 197134
rect 192576 162172 192628 162178
rect 192576 162114 192628 162120
rect 192760 148164 192812 148170
rect 192760 148106 192812 148112
rect 192666 141944 192722 141953
rect 192666 141879 192722 141888
rect 192574 140448 192630 140457
rect 192574 140383 192630 140392
rect 192484 76900 192536 76906
rect 192484 76842 192536 76848
rect 192588 72729 192616 140383
rect 192680 80578 192708 141879
rect 192772 138922 192800 148106
rect 192864 143585 192892 262482
rect 193128 197328 193180 197334
rect 193128 197270 193180 197276
rect 193140 197130 193168 197270
rect 193128 197124 193180 197130
rect 193128 197066 193180 197072
rect 193232 195974 193260 700334
rect 193864 547936 193916 547942
rect 193864 547878 193916 547884
rect 193876 265742 193904 547878
rect 193864 265736 193916 265742
rect 193864 265678 193916 265684
rect 193588 263628 193640 263634
rect 193588 263570 193640 263576
rect 193312 262472 193364 262478
rect 193312 262414 193364 262420
rect 193220 195968 193272 195974
rect 193220 195910 193272 195916
rect 192944 195900 192996 195906
rect 192944 195842 192996 195848
rect 192850 143576 192906 143585
rect 192850 143511 192906 143520
rect 192760 138916 192812 138922
rect 192760 138858 192812 138864
rect 192668 80572 192720 80578
rect 192668 80514 192720 80520
rect 192956 75818 192984 195842
rect 193220 189712 193272 189718
rect 193220 189654 193272 189660
rect 193128 182232 193180 182238
rect 193128 182174 193180 182180
rect 193140 182102 193168 182174
rect 193128 182096 193180 182102
rect 193128 182038 193180 182044
rect 192944 75812 192996 75818
rect 192944 75754 192996 75760
rect 192574 72720 192630 72729
rect 192574 72655 192630 72664
rect 192392 72412 192444 72418
rect 192392 72354 192444 72360
rect 192206 67008 192262 67017
rect 192206 66943 192262 66952
rect 192116 65952 192168 65958
rect 192116 65894 192168 65900
rect 193128 65952 193180 65958
rect 193128 65894 193180 65900
rect 193140 65686 193168 65894
rect 193128 65680 193180 65686
rect 193128 65622 193180 65628
rect 191288 64116 191340 64122
rect 191288 64058 191340 64064
rect 193232 62082 193260 189654
rect 193324 142118 193352 262414
rect 193404 262268 193456 262274
rect 193404 262210 193456 262216
rect 193416 143018 193444 262210
rect 193496 260908 193548 260914
rect 193496 260850 193548 260856
rect 193508 143138 193536 260850
rect 193600 145790 193628 263570
rect 193772 260296 193824 260302
rect 193772 260238 193824 260244
rect 193680 190188 193732 190194
rect 193680 190130 193732 190136
rect 193588 145784 193640 145790
rect 193588 145726 193640 145732
rect 193496 143132 193548 143138
rect 193496 143074 193548 143080
rect 193416 142990 193628 143018
rect 193600 142497 193628 142990
rect 193586 142488 193642 142497
rect 193586 142423 193642 142432
rect 193312 142112 193364 142118
rect 193312 142054 193364 142060
rect 193324 141438 193352 142054
rect 193404 141976 193456 141982
rect 193404 141918 193456 141924
rect 193312 141432 193364 141438
rect 193312 141374 193364 141380
rect 193416 70378 193444 141918
rect 193496 140344 193548 140350
rect 193496 140286 193548 140292
rect 193404 70372 193456 70378
rect 193404 70314 193456 70320
rect 193508 68678 193536 140286
rect 193600 140078 193628 142423
rect 193588 140072 193640 140078
rect 193588 140014 193640 140020
rect 193588 139936 193640 139942
rect 193588 139878 193640 139884
rect 193600 74050 193628 139878
rect 193588 74044 193640 74050
rect 193588 73986 193640 73992
rect 193692 73166 193720 190130
rect 193784 143002 193812 260238
rect 194520 200326 194548 700402
rect 194612 262886 194640 703582
rect 195624 703474 195652 703582
rect 195766 703520 195878 704960
rect 199630 703520 199742 704960
rect 202892 703582 203380 703610
rect 195808 703474 195836 703520
rect 195624 703446 195836 703474
rect 195980 700664 196032 700670
rect 195980 700606 196032 700612
rect 194692 700528 194744 700534
rect 194692 700470 194744 700476
rect 194600 262880 194652 262886
rect 194600 262822 194652 262828
rect 194508 200320 194560 200326
rect 194508 200262 194560 200268
rect 194520 198558 194548 200262
rect 194508 198552 194560 198558
rect 194508 198494 194560 198500
rect 194598 195392 194654 195401
rect 194598 195327 194654 195336
rect 193956 191276 194008 191282
rect 193956 191218 194008 191224
rect 193864 187264 193916 187270
rect 193864 187206 193916 187212
rect 193772 142996 193824 143002
rect 193772 142938 193824 142944
rect 193772 141772 193824 141778
rect 193772 141714 193824 141720
rect 193680 73160 193732 73166
rect 193680 73102 193732 73108
rect 193496 68672 193548 68678
rect 193496 68614 193548 68620
rect 193784 68474 193812 141714
rect 193876 74118 193904 187206
rect 193968 80889 193996 191218
rect 194048 147212 194100 147218
rect 194048 147154 194100 147160
rect 194060 105466 194088 147154
rect 194232 144356 194284 144362
rect 194232 144298 194284 144304
rect 194048 105460 194100 105466
rect 194048 105402 194100 105408
rect 194244 81122 194272 144298
rect 194232 81116 194284 81122
rect 194232 81058 194284 81064
rect 193954 80880 194010 80889
rect 193954 80815 194010 80824
rect 193864 74112 193916 74118
rect 193864 74054 193916 74060
rect 194612 72554 194640 195327
rect 194704 192846 194732 700470
rect 195244 276684 195296 276690
rect 195244 276626 195296 276632
rect 195256 276078 195284 276626
rect 195244 276072 195296 276078
rect 195244 276014 195296 276020
rect 195256 267734 195284 276014
rect 195256 267706 195376 267734
rect 194968 260364 195020 260370
rect 194968 260306 195020 260312
rect 194692 192840 194744 192846
rect 194692 192782 194744 192788
rect 194876 190256 194928 190262
rect 194876 190198 194928 190204
rect 194888 189854 194916 190198
rect 194876 189848 194928 189854
rect 194876 189790 194928 189796
rect 194888 180794 194916 189790
rect 194704 180766 194916 180794
rect 194704 72894 194732 180766
rect 194784 148980 194836 148986
rect 194784 148922 194836 148928
rect 194692 72888 194744 72894
rect 194692 72830 194744 72836
rect 194600 72548 194652 72554
rect 194600 72490 194652 72496
rect 193772 68468 193824 68474
rect 193772 68410 193824 68416
rect 194796 67318 194824 148922
rect 194876 144492 194928 144498
rect 194876 144434 194928 144440
rect 194888 68814 194916 144434
rect 194980 143070 195008 260306
rect 195244 259616 195296 259622
rect 195244 259558 195296 259564
rect 195060 259480 195112 259486
rect 195060 259422 195112 259428
rect 195072 143274 195100 259422
rect 195152 190052 195204 190058
rect 195152 189994 195204 190000
rect 195060 143268 195112 143274
rect 195060 143210 195112 143216
rect 194968 143064 195020 143070
rect 194968 143006 195020 143012
rect 195164 75546 195192 189994
rect 195256 145654 195284 259558
rect 195348 145897 195376 267706
rect 195426 259584 195482 259593
rect 195426 259519 195482 259528
rect 195334 145888 195390 145897
rect 195334 145823 195390 145832
rect 195244 145648 195296 145654
rect 195244 145590 195296 145596
rect 195440 142633 195468 259519
rect 195992 198626 196020 700606
rect 199384 700392 199436 700398
rect 199384 700334 199436 700340
rect 196624 648644 196676 648650
rect 196624 648586 196676 648592
rect 196636 263673 196664 648586
rect 198004 592068 198056 592074
rect 198004 592010 198056 592016
rect 198016 266694 198044 592010
rect 196992 266688 197044 266694
rect 196992 266630 197044 266636
rect 198004 266688 198056 266694
rect 198004 266630 198056 266636
rect 197004 266422 197032 266630
rect 198740 266484 198792 266490
rect 198740 266426 198792 266432
rect 196992 266416 197044 266422
rect 196992 266358 197044 266364
rect 196622 263664 196678 263673
rect 196622 263599 196678 263608
rect 196256 263016 196308 263022
rect 196256 262958 196308 262964
rect 196268 262342 196296 262958
rect 196256 262336 196308 262342
rect 196256 262278 196308 262284
rect 195980 198620 196032 198626
rect 195980 198562 196032 198568
rect 195992 194342 196020 198562
rect 195980 194336 196032 194342
rect 195980 194278 196032 194284
rect 195980 193928 196032 193934
rect 195980 193870 196032 193876
rect 195520 144560 195572 144566
rect 195520 144502 195572 144508
rect 195426 142624 195482 142633
rect 195426 142559 195482 142568
rect 195336 140548 195388 140554
rect 195336 140490 195388 140496
rect 195242 139224 195298 139233
rect 195242 139159 195298 139168
rect 195256 78198 195284 139159
rect 195348 80782 195376 140490
rect 195426 137456 195482 137465
rect 195426 137391 195482 137400
rect 195336 80776 195388 80782
rect 195336 80718 195388 80724
rect 195440 78305 195468 137391
rect 195426 78296 195482 78305
rect 195426 78231 195482 78240
rect 195244 78192 195296 78198
rect 195244 78134 195296 78140
rect 195152 75540 195204 75546
rect 195152 75482 195204 75488
rect 194876 68808 194928 68814
rect 194876 68750 194928 68756
rect 195532 68610 195560 144502
rect 195612 144424 195664 144430
rect 195612 144366 195664 144372
rect 195624 77926 195652 144366
rect 195612 77920 195664 77926
rect 195612 77862 195664 77868
rect 195992 72826 196020 193870
rect 196164 191344 196216 191350
rect 196164 191286 196216 191292
rect 196072 147280 196124 147286
rect 196072 147222 196124 147228
rect 195980 72820 196032 72826
rect 195980 72762 196032 72768
rect 195520 68604 195572 68610
rect 195520 68546 195572 68552
rect 194784 67312 194836 67318
rect 194784 67254 194836 67260
rect 196084 64462 196112 147222
rect 196176 74186 196204 191286
rect 196268 145450 196296 262278
rect 196440 260024 196492 260030
rect 196440 259966 196492 259972
rect 196256 145444 196308 145450
rect 196256 145386 196308 145392
rect 196452 145382 196480 259966
rect 196624 193996 196676 194002
rect 196624 193938 196676 193944
rect 196532 186992 196584 186998
rect 196532 186934 196584 186940
rect 196440 145376 196492 145382
rect 196440 145318 196492 145324
rect 196348 144900 196400 144906
rect 196348 144842 196400 144848
rect 196256 144764 196308 144770
rect 196256 144706 196308 144712
rect 196268 144226 196296 144706
rect 196256 144220 196308 144226
rect 196256 144162 196308 144168
rect 196164 74180 196216 74186
rect 196164 74122 196216 74128
rect 196360 70990 196388 144842
rect 196440 138780 196492 138786
rect 196440 138722 196492 138728
rect 196348 70984 196400 70990
rect 196348 70926 196400 70932
rect 196452 68882 196480 138722
rect 196544 74390 196572 186934
rect 196636 124914 196664 193938
rect 196900 148708 196952 148714
rect 196900 148650 196952 148656
rect 196808 145580 196860 145586
rect 196808 145522 196860 145528
rect 196716 140616 196768 140622
rect 196716 140558 196768 140564
rect 196624 124908 196676 124914
rect 196624 124850 196676 124856
rect 196532 74384 196584 74390
rect 196532 74326 196584 74332
rect 196728 73030 196756 140558
rect 196820 78130 196848 145522
rect 196808 78124 196860 78130
rect 196808 78066 196860 78072
rect 196716 73024 196768 73030
rect 196716 72966 196768 72972
rect 196440 68876 196492 68882
rect 196440 68818 196492 68824
rect 196912 68542 196940 148650
rect 197004 145625 197032 266358
rect 197360 265872 197412 265878
rect 197360 265814 197412 265820
rect 197084 259684 197136 259690
rect 197084 259626 197136 259632
rect 196990 145616 197046 145625
rect 196990 145551 197046 145560
rect 197096 144226 197124 259626
rect 197372 197985 197400 265814
rect 197636 262880 197688 262886
rect 197636 262822 197688 262828
rect 197544 262676 197596 262682
rect 197544 262618 197596 262624
rect 197358 197976 197414 197985
rect 197358 197911 197414 197920
rect 197452 195968 197504 195974
rect 197452 195910 197504 195916
rect 197360 192500 197412 192506
rect 197360 192442 197412 192448
rect 197084 144220 197136 144226
rect 197084 144162 197136 144168
rect 196900 68536 196952 68542
rect 196900 68478 196952 68484
rect 196072 64456 196124 64462
rect 196072 64398 196124 64404
rect 193220 62076 193272 62082
rect 193220 62018 193272 62024
rect 194508 62076 194560 62082
rect 194508 62018 194560 62024
rect 194520 61402 194548 62018
rect 194508 61396 194560 61402
rect 194508 61338 194560 61344
rect 190644 48272 190696 48278
rect 190644 48214 190696 48220
rect 191748 48272 191800 48278
rect 191748 48214 191800 48220
rect 191760 47666 191788 48214
rect 191748 47660 191800 47666
rect 191748 47602 191800 47608
rect 193220 40724 193272 40730
rect 193220 40666 193272 40672
rect 193232 16574 193260 40666
rect 197372 37262 197400 192442
rect 197464 74254 197492 195910
rect 197556 145602 197584 262618
rect 197648 145722 197676 262822
rect 197728 259956 197780 259962
rect 197728 259898 197780 259904
rect 197636 145716 197688 145722
rect 197636 145658 197688 145664
rect 197556 145574 197676 145602
rect 197544 144900 197596 144906
rect 197544 144842 197596 144848
rect 197556 144090 197584 144842
rect 197544 144084 197596 144090
rect 197544 144026 197596 144032
rect 197648 143206 197676 145574
rect 197740 144906 197768 259898
rect 197912 259888 197964 259894
rect 197912 259830 197964 259836
rect 197820 259752 197872 259758
rect 197820 259694 197872 259700
rect 197832 146062 197860 259694
rect 197924 146266 197952 259830
rect 198004 187332 198056 187338
rect 198004 187274 198056 187280
rect 197912 146260 197964 146266
rect 197912 146202 197964 146208
rect 197820 146056 197872 146062
rect 197820 145998 197872 146004
rect 197728 144900 197780 144906
rect 197728 144842 197780 144848
rect 197636 143200 197688 143206
rect 197636 143142 197688 143148
rect 197910 140720 197966 140729
rect 197910 140655 197966 140664
rect 197820 140412 197872 140418
rect 197820 140354 197872 140360
rect 197726 139088 197782 139097
rect 197726 139023 197782 139032
rect 197544 137828 197596 137834
rect 197544 137770 197596 137776
rect 197452 74248 197504 74254
rect 197452 74190 197504 74196
rect 197556 55214 197584 137770
rect 197740 67114 197768 139023
rect 197832 69630 197860 140354
rect 197924 71466 197952 140655
rect 198016 79354 198044 187274
rect 198096 153876 198148 153882
rect 198096 153818 198148 153824
rect 198108 153270 198136 153818
rect 198096 153264 198148 153270
rect 198096 153206 198148 153212
rect 198004 79348 198056 79354
rect 198004 79290 198056 79296
rect 197912 71460 197964 71466
rect 197912 71402 197964 71408
rect 197820 69624 197872 69630
rect 197820 69566 197872 69572
rect 198108 67454 198136 153206
rect 198280 148844 198332 148850
rect 198280 148786 198332 148792
rect 198188 144152 198240 144158
rect 198188 144094 198240 144100
rect 198200 91118 198228 144094
rect 198188 91112 198240 91118
rect 198188 91054 198240 91060
rect 198096 67448 198148 67454
rect 198096 67390 198148 67396
rect 197728 67108 197780 67114
rect 197728 67050 197780 67056
rect 198292 55214 198320 148786
rect 198752 145926 198780 266426
rect 198924 263696 198976 263702
rect 198924 263638 198976 263644
rect 198830 196480 198886 196489
rect 198830 196415 198886 196424
rect 198844 195770 198872 196415
rect 198832 195764 198884 195770
rect 198832 195706 198884 195712
rect 198832 193996 198884 194002
rect 198832 193938 198884 193944
rect 198844 192953 198872 193938
rect 198830 192944 198886 192953
rect 198830 192879 198886 192888
rect 198740 145920 198792 145926
rect 198740 145862 198792 145868
rect 198844 72593 198872 192879
rect 198936 145858 198964 263638
rect 199108 262608 199160 262614
rect 199108 262550 199160 262556
rect 199016 184476 199068 184482
rect 199016 184418 199068 184424
rect 198924 145852 198976 145858
rect 198924 145794 198976 145800
rect 198830 72584 198886 72593
rect 198830 72519 198886 72528
rect 199028 67250 199056 184418
rect 199120 146130 199148 262550
rect 199396 199578 199424 700334
rect 199672 699718 199700 703520
rect 200120 700596 200172 700602
rect 200120 700538 200172 700544
rect 199660 699712 199712 699718
rect 199660 699654 199712 699660
rect 199384 199572 199436 199578
rect 199384 199514 199436 199520
rect 199200 190528 199252 190534
rect 199200 190470 199252 190476
rect 199108 146124 199160 146130
rect 199108 146066 199160 146072
rect 199108 140480 199160 140486
rect 199108 140422 199160 140428
rect 199016 67244 199068 67250
rect 199016 67186 199068 67192
rect 199120 67182 199148 140422
rect 199212 75041 199240 190470
rect 199384 187672 199436 187678
rect 199384 187614 199436 187620
rect 199292 184408 199344 184414
rect 199292 184350 199344 184356
rect 199198 75032 199254 75041
rect 199198 74967 199254 74976
rect 199304 73982 199332 184350
rect 199396 81297 199424 187614
rect 200132 187513 200160 700538
rect 201500 699712 201552 699718
rect 201500 699654 201552 699660
rect 200764 560312 200816 560318
rect 200764 560254 200816 560260
rect 200776 269822 200804 560254
rect 200764 269816 200816 269822
rect 200764 269758 200816 269764
rect 201408 199504 201460 199510
rect 201408 199446 201460 199452
rect 201420 198694 201448 199446
rect 200396 198688 200448 198694
rect 200396 198630 200448 198636
rect 201408 198688 201460 198694
rect 201408 198630 201460 198636
rect 200212 197056 200264 197062
rect 200212 196998 200264 197004
rect 200118 187504 200174 187513
rect 200118 187439 200174 187448
rect 199660 148912 199712 148918
rect 199660 148854 199712 148860
rect 199568 144832 199620 144838
rect 199568 144774 199620 144780
rect 199474 138680 199530 138689
rect 199474 138615 199530 138624
rect 199382 81288 199438 81297
rect 199382 81223 199438 81232
rect 199292 73976 199344 73982
rect 199292 73918 199344 73924
rect 199108 67176 199160 67182
rect 199108 67118 199160 67124
rect 199488 65657 199516 138615
rect 199580 71058 199608 144774
rect 199568 71052 199620 71058
rect 199568 70994 199620 71000
rect 199672 68406 199700 148854
rect 199752 146192 199804 146198
rect 199752 146134 199804 146140
rect 199764 71194 199792 146134
rect 199752 71188 199804 71194
rect 199752 71130 199804 71136
rect 200224 70174 200252 196998
rect 200304 195628 200356 195634
rect 200304 195570 200356 195576
rect 200316 187678 200344 195570
rect 200304 187672 200356 187678
rect 200304 187614 200356 187620
rect 200408 76537 200436 198630
rect 200488 194132 200540 194138
rect 200488 194074 200540 194080
rect 200500 77246 200528 194074
rect 201512 192982 201540 699654
rect 202144 665236 202196 665242
rect 202144 665178 202196 665184
rect 202156 271250 202184 665178
rect 202144 271244 202196 271250
rect 202144 271186 202196 271192
rect 202236 194676 202288 194682
rect 202236 194618 202288 194624
rect 202248 194177 202276 194618
rect 202234 194168 202290 194177
rect 202234 194103 202290 194112
rect 201500 192976 201552 192982
rect 201500 192918 201552 192924
rect 201590 192808 201646 192817
rect 201590 192743 201646 192752
rect 200856 191548 200908 191554
rect 200856 191490 200908 191496
rect 200580 187400 200632 187406
rect 200580 187342 200632 187348
rect 200488 77240 200540 77246
rect 200488 77182 200540 77188
rect 200394 76528 200450 76537
rect 200394 76463 200450 76472
rect 200592 73953 200620 187342
rect 200672 148300 200724 148306
rect 200672 148242 200724 148248
rect 200578 73944 200634 73953
rect 200578 73879 200634 73888
rect 200212 70168 200264 70174
rect 200212 70110 200264 70116
rect 199660 68400 199712 68406
rect 199660 68342 199712 68348
rect 200210 67008 200266 67017
rect 200210 66943 200212 66952
rect 200264 66943 200266 66952
rect 200212 66914 200264 66920
rect 200684 65754 200712 148242
rect 200762 137320 200818 137329
rect 200762 137255 200818 137264
rect 200672 65748 200724 65754
rect 200672 65690 200724 65696
rect 199474 65648 199530 65657
rect 199474 65583 199530 65592
rect 200776 64705 200804 137255
rect 200868 137154 200896 191490
rect 201038 191312 201094 191321
rect 201038 191247 201094 191256
rect 200948 146328 201000 146334
rect 200948 146270 201000 146276
rect 200856 137148 200908 137154
rect 200856 137090 200908 137096
rect 200854 134464 200910 134473
rect 200854 134399 200910 134408
rect 200868 64734 200896 134399
rect 200960 81841 200988 146270
rect 200946 81832 201002 81841
rect 200946 81767 201002 81776
rect 201052 67289 201080 191247
rect 201132 187604 201184 187610
rect 201132 187546 201184 187552
rect 201038 67280 201094 67289
rect 201038 67215 201094 67224
rect 200856 64728 200908 64734
rect 200762 64696 200818 64705
rect 200856 64670 200908 64676
rect 200762 64631 200818 64640
rect 201144 59294 201172 187546
rect 201408 187400 201460 187406
rect 201408 187342 201460 187348
rect 201420 186998 201448 187342
rect 201498 187096 201554 187105
rect 201498 187031 201554 187040
rect 201408 186992 201460 186998
rect 201408 186934 201460 186940
rect 201408 147144 201460 147150
rect 201408 147086 201460 147092
rect 201420 146334 201448 147086
rect 201408 146328 201460 146334
rect 201408 146270 201460 146276
rect 201512 71505 201540 187031
rect 201498 71496 201554 71505
rect 201498 71431 201554 71440
rect 201498 70272 201554 70281
rect 201498 70207 201554 70216
rect 201512 69970 201540 70207
rect 201500 69964 201552 69970
rect 201500 69906 201552 69912
rect 201604 67153 201632 192743
rect 201776 187536 201828 187542
rect 201776 187478 201828 187484
rect 201684 187468 201736 187474
rect 201684 187410 201736 187416
rect 201696 73642 201724 187410
rect 201788 75410 201816 187478
rect 202892 183394 202920 703582
rect 203352 703474 203380 703582
rect 203494 703520 203606 704960
rect 207032 703582 207244 703610
rect 203536 703474 203564 703520
rect 203352 703446 203564 703474
rect 206284 350600 206336 350606
rect 206284 350542 206336 350548
rect 206296 272542 206324 350542
rect 206284 272536 206336 272542
rect 206284 272478 206336 272484
rect 204260 201544 204312 201550
rect 204260 201486 204312 201492
rect 202972 194472 203024 194478
rect 202972 194414 203024 194420
rect 202880 183388 202932 183394
rect 202880 183330 202932 183336
rect 201868 178832 201920 178838
rect 201868 178774 201920 178780
rect 201880 79422 201908 178774
rect 201960 148776 202012 148782
rect 201960 148718 202012 148724
rect 201868 79416 201920 79422
rect 201868 79358 201920 79364
rect 201776 75404 201828 75410
rect 201776 75346 201828 75352
rect 201684 73636 201736 73642
rect 201684 73578 201736 73584
rect 201684 71256 201736 71262
rect 201684 71198 201736 71204
rect 201590 67144 201646 67153
rect 201590 67079 201646 67088
rect 201696 64874 201724 71198
rect 201972 65618 202000 148718
rect 202052 148640 202104 148646
rect 202052 148582 202104 148588
rect 202064 68134 202092 148582
rect 202144 148232 202196 148238
rect 202144 148174 202196 148180
rect 202156 71262 202184 148174
rect 202236 138916 202288 138922
rect 202236 138858 202288 138864
rect 202144 71256 202196 71262
rect 202144 71198 202196 71204
rect 202052 68128 202104 68134
rect 202052 68070 202104 68076
rect 201960 65612 202012 65618
rect 201960 65554 202012 65560
rect 201512 64846 201724 64874
rect 201132 59288 201184 59294
rect 201132 59230 201184 59236
rect 201408 59288 201460 59294
rect 201408 59230 201460 59236
rect 201420 58750 201448 59230
rect 201408 58744 201460 58750
rect 201408 58686 201460 58692
rect 197464 55186 197584 55214
rect 198280 55208 198332 55214
rect 197464 51066 197492 55186
rect 198280 55150 198332 55156
rect 198292 54534 198320 55150
rect 198280 54528 198332 54534
rect 198280 54470 198332 54476
rect 197452 51060 197504 51066
rect 197452 51002 197504 51008
rect 197464 50386 197492 51002
rect 197452 50380 197504 50386
rect 197452 50322 197504 50328
rect 197360 37256 197412 37262
rect 197360 37198 197412 37204
rect 201512 16574 201540 64846
rect 202248 62762 202276 138858
rect 202328 105460 202380 105466
rect 202328 105402 202380 105408
rect 202340 80034 202368 105402
rect 202878 81152 202934 81161
rect 202878 81087 202934 81096
rect 202892 81054 202920 81087
rect 202880 81048 202932 81054
rect 202880 80990 202932 80996
rect 202328 80028 202380 80034
rect 202328 79970 202380 79976
rect 202788 80028 202840 80034
rect 202788 79970 202840 79976
rect 202800 79082 202828 79970
rect 202788 79076 202840 79082
rect 202788 79018 202840 79024
rect 202788 75404 202840 75410
rect 202788 75346 202840 75352
rect 202800 75274 202828 75346
rect 202788 75268 202840 75274
rect 202788 75210 202840 75216
rect 202984 73778 203012 194414
rect 203064 194064 203116 194070
rect 203064 194006 203116 194012
rect 203076 76634 203104 194006
rect 203432 188284 203484 188290
rect 203432 188226 203484 188232
rect 203156 187196 203208 187202
rect 203156 187138 203208 187144
rect 203064 76628 203116 76634
rect 203064 76570 203116 76576
rect 202972 73772 203024 73778
rect 202972 73714 203024 73720
rect 203168 71330 203196 187138
rect 203340 185972 203392 185978
rect 203340 185914 203392 185920
rect 203248 178900 203300 178906
rect 203248 178842 203300 178848
rect 203156 71324 203208 71330
rect 203156 71266 203208 71272
rect 203260 66026 203288 178842
rect 203352 76702 203380 185914
rect 203444 81025 203472 188226
rect 203892 184680 203944 184686
rect 203892 184622 203944 184628
rect 203616 148572 203668 148578
rect 203616 148514 203668 148520
rect 203522 148472 203578 148481
rect 203522 148407 203578 148416
rect 203430 81016 203486 81025
rect 203430 80951 203486 80960
rect 203340 76696 203392 76702
rect 203340 76638 203392 76644
rect 203248 66020 203300 66026
rect 203248 65962 203300 65968
rect 202236 62756 202288 62762
rect 202236 62698 202288 62704
rect 203536 59362 203564 148407
rect 203628 68270 203656 148514
rect 203708 137148 203760 137154
rect 203708 137090 203760 137096
rect 203720 136678 203748 137090
rect 203708 136672 203760 136678
rect 203708 136614 203760 136620
rect 203720 80986 203748 136614
rect 203708 80980 203760 80986
rect 203708 80922 203760 80928
rect 203800 80096 203852 80102
rect 203800 80038 203852 80044
rect 203812 73098 203840 80038
rect 203800 73092 203852 73098
rect 203800 73034 203852 73040
rect 203616 68264 203668 68270
rect 203616 68206 203668 68212
rect 203904 64394 203932 184622
rect 204272 71534 204300 201486
rect 204352 200864 204404 200870
rect 204352 200806 204404 200812
rect 204364 200190 204392 200806
rect 204352 200184 204404 200190
rect 204352 200126 204404 200132
rect 204260 71528 204312 71534
rect 204260 71470 204312 71476
rect 204258 70272 204314 70281
rect 204258 70207 204314 70216
rect 204272 69902 204300 70207
rect 204364 70009 204392 200126
rect 207032 194410 207060 703582
rect 207216 703474 207244 703582
rect 207358 703520 207470 704960
rect 211222 703520 211334 704960
rect 213932 703582 214972 703610
rect 207400 703474 207428 703520
rect 207216 703446 207428 703474
rect 210424 415472 210476 415478
rect 210424 415414 210476 415420
rect 210436 266014 210464 415414
rect 210424 266008 210476 266014
rect 210424 265950 210476 265956
rect 211436 200320 211488 200326
rect 211436 200262 211488 200268
rect 208400 198212 208452 198218
rect 208400 198154 208452 198160
rect 207112 196648 207164 196654
rect 207112 196590 207164 196596
rect 207020 194404 207072 194410
rect 207020 194346 207072 194352
rect 204444 194336 204496 194342
rect 204444 194278 204496 194284
rect 204456 72622 204484 194278
rect 205640 194200 205692 194206
rect 205640 194142 205692 194148
rect 204720 192840 204772 192846
rect 204720 192782 204772 192788
rect 204536 184748 204588 184754
rect 204536 184690 204588 184696
rect 204444 72616 204496 72622
rect 204444 72558 204496 72564
rect 204350 70000 204406 70009
rect 204350 69935 204406 69944
rect 204260 69896 204312 69902
rect 204260 69838 204312 69844
rect 204548 67046 204576 184690
rect 204628 184544 204680 184550
rect 204628 184486 204680 184492
rect 204640 68377 204668 184486
rect 204732 80102 204760 192782
rect 204812 184068 204864 184074
rect 204812 184010 204864 184016
rect 204720 80096 204772 80102
rect 204720 80038 204772 80044
rect 204824 76430 204852 184010
rect 204996 148504 205048 148510
rect 204996 148446 205048 148452
rect 204904 140208 204956 140214
rect 204904 140150 204956 140156
rect 204812 76424 204864 76430
rect 204812 76366 204864 76372
rect 204626 68368 204682 68377
rect 204626 68303 204682 68312
rect 204536 67040 204588 67046
rect 204536 66982 204588 66988
rect 203892 64388 203944 64394
rect 203892 64330 203944 64336
rect 203524 59356 203576 59362
rect 203524 59298 203576 59304
rect 204168 59356 204220 59362
rect 204168 59298 204220 59304
rect 204180 58682 204208 59298
rect 204168 58676 204220 58682
rect 204168 58618 204220 58624
rect 204916 57934 204944 140150
rect 205008 78062 205036 148446
rect 205088 138848 205140 138854
rect 205088 138790 205140 138796
rect 205100 81705 205128 138790
rect 205086 81696 205142 81705
rect 205086 81631 205142 81640
rect 204996 78056 205048 78062
rect 204996 77998 205048 78004
rect 205652 70106 205680 194142
rect 206468 189100 206520 189106
rect 206468 189042 206520 189048
rect 205824 188692 205876 188698
rect 205824 188634 205876 188640
rect 205732 184612 205784 184618
rect 205732 184554 205784 184560
rect 205640 70100 205692 70106
rect 205640 70042 205692 70048
rect 205638 70000 205694 70009
rect 205638 69935 205694 69944
rect 205652 69834 205680 69935
rect 205640 69828 205692 69834
rect 205640 69770 205692 69776
rect 205744 64802 205772 184554
rect 205836 68921 205864 188634
rect 206480 188562 206508 189042
rect 206008 188556 206060 188562
rect 206008 188498 206060 188504
rect 206468 188556 206520 188562
rect 206468 188498 206520 188504
rect 205916 181960 205968 181966
rect 205916 181902 205968 181908
rect 205822 68912 205878 68921
rect 205822 68847 205878 68856
rect 205732 64796 205784 64802
rect 205732 64738 205784 64744
rect 205928 64598 205956 181902
rect 206020 71602 206048 188498
rect 207020 185836 207072 185842
rect 207020 185778 207072 185784
rect 206100 184340 206152 184346
rect 206100 184282 206152 184288
rect 206008 71596 206060 71602
rect 206008 71538 206060 71544
rect 206112 68241 206140 184282
rect 206192 162172 206244 162178
rect 206192 162114 206244 162120
rect 206204 161498 206232 162114
rect 206192 161492 206244 161498
rect 206192 161434 206244 161440
rect 206204 78470 206232 161434
rect 206376 147076 206428 147082
rect 206376 147018 206428 147024
rect 206284 141568 206336 141574
rect 206284 141510 206336 141516
rect 206192 78464 206244 78470
rect 206192 78406 206244 78412
rect 206098 68232 206154 68241
rect 206098 68167 206154 68176
rect 205916 64592 205968 64598
rect 205916 64534 205968 64540
rect 206296 63102 206324 141510
rect 206388 77994 206416 147018
rect 206468 124908 206520 124914
rect 206468 124850 206520 124856
rect 206480 124234 206508 124850
rect 206468 124228 206520 124234
rect 206468 124170 206520 124176
rect 206480 82142 206508 124170
rect 206468 82136 206520 82142
rect 206468 82078 206520 82084
rect 206376 77988 206428 77994
rect 206376 77930 206428 77936
rect 207032 64530 207060 185778
rect 207124 71602 207152 196590
rect 207296 195696 207348 195702
rect 207296 195638 207348 195644
rect 207204 183184 207256 183190
rect 207204 183126 207256 183132
rect 207112 71596 207164 71602
rect 207112 71538 207164 71544
rect 207110 71496 207166 71505
rect 207110 71431 207166 71440
rect 207124 71398 207152 71431
rect 207112 71392 207164 71398
rect 207112 71334 207164 71340
rect 207020 64524 207072 64530
rect 207020 64466 207072 64472
rect 206284 63096 206336 63102
rect 206284 63038 206336 63044
rect 207216 62966 207244 183126
rect 207308 75138 207336 195638
rect 208412 192930 208440 198154
rect 209872 197260 209924 197266
rect 209872 197202 209924 197208
rect 208492 196988 208544 196994
rect 208492 196930 208544 196936
rect 208320 192902 208440 192930
rect 208320 192386 208348 192902
rect 208400 192772 208452 192778
rect 208400 192714 208452 192720
rect 208412 192506 208440 192714
rect 208400 192500 208452 192506
rect 208400 192442 208452 192448
rect 208320 192358 208440 192386
rect 207388 188624 207440 188630
rect 207388 188566 207440 188572
rect 207400 80918 207428 188566
rect 207478 187232 207534 187241
rect 207478 187167 207534 187176
rect 207492 81297 207520 187167
rect 207664 149048 207716 149054
rect 207664 148990 207716 148996
rect 207572 144220 207624 144226
rect 207572 144162 207624 144168
rect 207478 81288 207534 81297
rect 207478 81223 207534 81232
rect 207388 80912 207440 80918
rect 207388 80854 207440 80860
rect 207296 75132 207348 75138
rect 207296 75074 207348 75080
rect 207296 71596 207348 71602
rect 207296 71538 207348 71544
rect 207308 69698 207336 71538
rect 207388 70032 207440 70038
rect 207388 69974 207440 69980
rect 207400 69698 207428 69974
rect 207296 69692 207348 69698
rect 207296 69634 207348 69640
rect 207388 69692 207440 69698
rect 207388 69634 207440 69640
rect 207584 64326 207612 144162
rect 207676 70038 207704 148990
rect 207848 142520 207900 142526
rect 207848 142462 207900 142468
rect 207754 141808 207810 141817
rect 207754 141743 207810 141752
rect 207768 70310 207796 141743
rect 207860 78538 207888 142462
rect 207848 78532 207900 78538
rect 207848 78474 207900 78480
rect 207756 70304 207808 70310
rect 207756 70246 207808 70252
rect 207664 70032 207716 70038
rect 207664 69974 207716 69980
rect 208412 65890 208440 192358
rect 208504 75614 208532 196930
rect 208584 195424 208636 195430
rect 208584 195366 208636 195372
rect 208492 75608 208544 75614
rect 208492 75550 208544 75556
rect 208596 75478 208624 195366
rect 209780 195288 209832 195294
rect 209780 195230 209832 195236
rect 208952 192500 209004 192506
rect 208952 192442 209004 192448
rect 208674 185736 208730 185745
rect 208674 185671 208730 185680
rect 208584 75472 208636 75478
rect 208584 75414 208636 75420
rect 208688 67386 208716 185671
rect 208768 181416 208820 181422
rect 208768 181358 208820 181364
rect 208676 67380 208728 67386
rect 208676 67322 208728 67328
rect 208400 65884 208452 65890
rect 208400 65826 208452 65832
rect 208780 64666 208808 181358
rect 208860 180192 208912 180198
rect 208860 180134 208912 180140
rect 208768 64660 208820 64666
rect 208768 64602 208820 64608
rect 207572 64320 207624 64326
rect 207572 64262 207624 64268
rect 208872 63034 208900 180134
rect 208964 76838 208992 192442
rect 209136 191208 209188 191214
rect 209136 191150 209188 191156
rect 209042 188592 209098 188601
rect 209042 188527 209098 188536
rect 208952 76832 209004 76838
rect 208952 76774 209004 76780
rect 209056 75857 209084 188527
rect 209148 79558 209176 191150
rect 209228 189916 209280 189922
rect 209228 189858 209280 189864
rect 209136 79552 209188 79558
rect 209136 79494 209188 79500
rect 209240 79218 209268 189858
rect 209228 79212 209280 79218
rect 209228 79154 209280 79160
rect 209042 75848 209098 75857
rect 209042 75783 209098 75792
rect 209792 66094 209820 195230
rect 209884 68785 209912 197202
rect 209964 197124 210016 197130
rect 209964 197066 210016 197072
rect 209976 78606 210004 197066
rect 211158 194984 211214 194993
rect 211158 194919 211214 194928
rect 210240 186924 210292 186930
rect 210240 186866 210292 186872
rect 210148 184952 210200 184958
rect 210148 184894 210200 184900
rect 210056 178764 210108 178770
rect 210056 178706 210108 178712
rect 209964 78600 210016 78606
rect 209964 78542 210016 78548
rect 209962 76800 210018 76809
rect 209962 76735 209964 76744
rect 210016 76735 210018 76744
rect 209964 76706 210016 76712
rect 209870 68776 209926 68785
rect 209870 68711 209926 68720
rect 209780 66088 209832 66094
rect 209780 66030 209832 66036
rect 210068 63238 210096 178706
rect 210160 71738 210188 184894
rect 210252 75342 210280 186866
rect 210424 185020 210476 185026
rect 210424 184962 210476 184968
rect 210332 181348 210384 181354
rect 210332 181290 210384 181296
rect 210240 75336 210292 75342
rect 210344 75313 210372 181290
rect 210436 79286 210464 184962
rect 210608 151292 210660 151298
rect 210608 151234 210660 151240
rect 210516 147008 210568 147014
rect 210516 146950 210568 146956
rect 210424 79280 210476 79286
rect 210424 79222 210476 79228
rect 210240 75278 210292 75284
rect 210330 75304 210386 75313
rect 210330 75239 210386 75248
rect 210148 71732 210200 71738
rect 210148 71674 210200 71680
rect 210056 63232 210108 63238
rect 210056 63174 210108 63180
rect 210528 63170 210556 146950
rect 210620 112470 210648 151234
rect 210608 112464 210660 112470
rect 210608 112406 210660 112412
rect 210620 79150 210648 112406
rect 210608 79144 210660 79150
rect 210608 79086 210660 79092
rect 211172 66881 211200 194919
rect 211252 185768 211304 185774
rect 211252 185710 211304 185716
rect 211158 66872 211214 66881
rect 211158 66807 211214 66816
rect 211264 63209 211292 185710
rect 211344 185564 211396 185570
rect 211344 185506 211396 185512
rect 211356 63481 211384 185506
rect 211448 77761 211476 200262
rect 212724 196920 212776 196926
rect 212724 196862 212776 196868
rect 212632 196852 212684 196858
rect 212632 196794 212684 196800
rect 212446 195800 212502 195809
rect 212446 195735 212502 195744
rect 211526 195664 211582 195673
rect 211526 195599 211582 195608
rect 211540 78878 211568 195599
rect 212460 194993 212488 195735
rect 212540 195356 212592 195362
rect 212540 195298 212592 195304
rect 212446 194984 212502 194993
rect 212446 194919 212502 194928
rect 211804 187128 211856 187134
rect 211804 187070 211856 187076
rect 211712 185904 211764 185910
rect 211712 185846 211764 185852
rect 211620 181892 211672 181898
rect 211620 181834 211672 181840
rect 211528 78872 211580 78878
rect 211528 78814 211580 78820
rect 211434 77752 211490 77761
rect 211434 77687 211490 77696
rect 211632 67522 211660 181834
rect 211724 74458 211752 185846
rect 211816 77042 211844 187070
rect 212448 185768 212500 185774
rect 212448 185710 212500 185716
rect 212460 185570 212488 185710
rect 212448 185564 212500 185570
rect 212448 185506 212500 185512
rect 211988 148436 212040 148442
rect 211988 148378 212040 148384
rect 211896 148368 211948 148374
rect 211896 148310 211948 148316
rect 211908 77110 211936 148310
rect 212000 80714 212028 148378
rect 211988 80708 212040 80714
rect 211988 80650 212040 80656
rect 211896 77104 211948 77110
rect 211896 77046 211948 77052
rect 211804 77036 211856 77042
rect 211804 76978 211856 76984
rect 211712 74452 211764 74458
rect 211712 74394 211764 74400
rect 211804 68332 211856 68338
rect 211804 68274 211856 68280
rect 211620 67516 211672 67522
rect 211620 67458 211672 67464
rect 211342 63472 211398 63481
rect 211342 63407 211398 63416
rect 211250 63200 211306 63209
rect 210516 63164 210568 63170
rect 211250 63135 211306 63144
rect 210516 63106 210568 63112
rect 208860 63028 208912 63034
rect 208860 62970 208912 62976
rect 207204 62960 207256 62966
rect 207204 62902 207256 62908
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 204916 57322 204944 57870
rect 204904 57316 204956 57322
rect 204904 57258 204956 57264
rect 205640 53168 205692 53174
rect 205640 53110 205692 53116
rect 193232 16546 194088 16574
rect 201512 16546 201816 16574
rect 190614 354 190726 480
rect 190472 326 190726 354
rect 194060 354 194088 16546
rect 194478 354 194590 480
rect 194060 326 194590 354
rect 190614 -960 190726 326
rect 194478 -960 194590 326
rect 198342 -960 198454 480
rect 201788 354 201816 16546
rect 202206 354 202318 480
rect 201788 326 202318 354
rect 205652 354 205680 53110
rect 211816 3058 211844 68274
rect 212448 67516 212500 67522
rect 212448 67458 212500 67464
rect 212460 66978 212488 67458
rect 212448 66972 212500 66978
rect 212448 66914 212500 66920
rect 212552 64870 212580 195298
rect 212644 75585 212672 196794
rect 212736 78946 212764 196862
rect 212816 195764 212868 195770
rect 212816 195706 212868 195712
rect 213828 195764 213880 195770
rect 213828 195706 213880 195712
rect 212828 79393 212856 195706
rect 213840 195362 213868 195706
rect 213828 195356 213880 195362
rect 213828 195298 213880 195304
rect 213000 183388 213052 183394
rect 213000 183330 213052 183336
rect 212908 183320 212960 183326
rect 212908 183262 212960 183268
rect 212814 79384 212870 79393
rect 212814 79319 212870 79328
rect 212724 78940 212776 78946
rect 212724 78882 212776 78888
rect 212630 75576 212686 75585
rect 212630 75511 212686 75520
rect 212920 70242 212948 183262
rect 213012 77790 213040 183330
rect 213092 183252 213144 183258
rect 213092 183194 213144 183200
rect 213104 78577 213132 183194
rect 213932 182034 213960 703582
rect 214944 703474 214972 703582
rect 215086 703520 215198 704960
rect 218072 703582 218836 703610
rect 215128 703474 215156 703520
rect 214944 703446 215156 703474
rect 218072 273970 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 222814 703520 222926 704960
rect 226678 703520 226790 704960
rect 230542 703520 230654 704960
rect 233252 703582 234292 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 222856 699718 222884 703520
rect 226720 699718 226748 703520
rect 220084 699712 220136 699718
rect 220084 699654 220136 699660
rect 222844 699712 222896 699718
rect 222844 699654 222896 699660
rect 224224 699712 224276 699718
rect 224224 699654 224276 699660
rect 226708 699712 226760 699718
rect 226708 699654 226760 699660
rect 218060 273964 218112 273970
rect 218060 273906 218112 273912
rect 215392 200252 215444 200258
rect 215392 200194 215444 200200
rect 214656 196784 214708 196790
rect 214656 196726 214708 196732
rect 214380 195424 214432 195430
rect 214380 195366 214432 195372
rect 214392 194682 214420 195366
rect 214012 194676 214064 194682
rect 214012 194618 214064 194624
rect 214380 194676 214432 194682
rect 214380 194618 214432 194624
rect 213920 182028 213972 182034
rect 213920 181970 213972 181976
rect 213090 78568 213146 78577
rect 213090 78503 213146 78512
rect 213000 77784 213052 77790
rect 213000 77726 213052 77732
rect 214024 75721 214052 194618
rect 214102 192672 214158 192681
rect 214102 192607 214158 192616
rect 214010 75712 214066 75721
rect 214010 75647 214066 75656
rect 214116 75206 214144 192607
rect 214288 192568 214340 192574
rect 214288 192510 214340 192516
rect 214194 178936 214250 178945
rect 214194 178871 214250 178880
rect 214104 75200 214156 75206
rect 214104 75142 214156 75148
rect 212908 70236 212960 70242
rect 212908 70178 212960 70184
rect 212540 64864 212592 64870
rect 212540 64806 212592 64812
rect 214208 63345 214236 178871
rect 214300 79966 214328 192510
rect 214378 189816 214434 189825
rect 214378 189751 214434 189760
rect 214288 79960 214340 79966
rect 214288 79902 214340 79908
rect 214392 78985 214420 189751
rect 214562 187504 214618 187513
rect 214562 187439 214618 187448
rect 214576 186833 214604 187439
rect 214562 186824 214618 186833
rect 214562 186759 214618 186768
rect 214576 180794 214604 186759
rect 214484 180766 214604 180794
rect 214378 78976 214434 78985
rect 214378 78911 214434 78920
rect 214484 78849 214512 180766
rect 214564 151156 214616 151162
rect 214564 151098 214616 151104
rect 214470 78840 214526 78849
rect 214470 78775 214526 78784
rect 214194 63336 214250 63345
rect 214194 63271 214250 63280
rect 214576 56574 214604 151098
rect 214668 149734 214696 196726
rect 215300 196716 215352 196722
rect 215300 196658 215352 196664
rect 215312 196042 215340 196658
rect 215300 196036 215352 196042
rect 215300 195978 215352 195984
rect 215300 195560 215352 195566
rect 215300 195502 215352 195508
rect 214840 182844 214892 182850
rect 214840 182786 214892 182792
rect 214656 149728 214708 149734
rect 214656 149670 214708 149676
rect 214668 75070 214696 149670
rect 214748 140140 214800 140146
rect 214748 140082 214800 140088
rect 214760 139466 214788 140082
rect 214748 139460 214800 139466
rect 214748 139402 214800 139408
rect 214656 75064 214708 75070
rect 214656 75006 214708 75012
rect 214760 75002 214788 139402
rect 214748 74996 214800 75002
rect 214748 74938 214800 74944
rect 214852 65385 214880 182786
rect 215312 71670 215340 195502
rect 215404 76401 215432 200194
rect 216680 199572 216732 199578
rect 216680 199514 216732 199520
rect 216692 199238 216720 199514
rect 216680 199232 216732 199238
rect 216680 199174 216732 199180
rect 215576 196036 215628 196042
rect 215576 195978 215628 195984
rect 215484 195492 215536 195498
rect 215484 195434 215536 195440
rect 215390 76392 215446 76401
rect 215390 76327 215446 76336
rect 215392 75744 215444 75750
rect 215392 75686 215444 75692
rect 215404 75206 215432 75686
rect 215496 75682 215524 195434
rect 215588 77178 215616 195978
rect 216692 190454 216720 199174
rect 219532 198144 219584 198150
rect 219532 198086 219584 198092
rect 219440 198076 219492 198082
rect 219440 198018 219492 198024
rect 218058 195528 218114 195537
rect 218058 195463 218114 195472
rect 217140 192636 217192 192642
rect 217140 192578 217192 192584
rect 216692 190426 216812 190454
rect 215852 188488 215904 188494
rect 215852 188430 215904 188436
rect 215760 182912 215812 182918
rect 215760 182854 215812 182860
rect 215668 181756 215720 181762
rect 215668 181698 215720 181704
rect 215576 77172 215628 77178
rect 215576 77114 215628 77120
rect 215484 75676 215536 75682
rect 215484 75618 215536 75624
rect 215392 75200 215444 75206
rect 215392 75142 215444 75148
rect 215300 71664 215352 71670
rect 215300 71606 215352 71612
rect 215312 71058 215340 71606
rect 215300 71052 215352 71058
rect 215300 70994 215352 71000
rect 214838 65376 214894 65385
rect 214838 65311 214894 65320
rect 215680 63374 215708 181698
rect 215772 65929 215800 182854
rect 215864 75750 215892 188430
rect 215944 185632 215996 185638
rect 215944 185574 215996 185580
rect 215956 77897 215984 185574
rect 216680 182980 216732 182986
rect 216680 182922 216732 182928
rect 216036 151088 216088 151094
rect 216036 151030 216088 151036
rect 215942 77888 215998 77897
rect 215942 77823 215998 77832
rect 215852 75744 215904 75750
rect 215852 75686 215904 75692
rect 215758 65920 215814 65929
rect 215758 65855 215814 65864
rect 215668 63368 215720 63374
rect 215668 63310 215720 63316
rect 214564 56568 214616 56574
rect 214564 56510 214616 56516
rect 214576 55962 214604 56510
rect 214564 55956 214616 55962
rect 214564 55898 214616 55904
rect 216048 46918 216076 151030
rect 216126 148336 216182 148345
rect 216126 148271 216182 148280
rect 216140 69018 216168 148271
rect 216128 69012 216180 69018
rect 216128 68954 216180 68960
rect 216692 66162 216720 182922
rect 216784 81977 216812 190426
rect 217046 185872 217102 185881
rect 217046 185807 217102 185816
rect 216956 184204 217008 184210
rect 216956 184146 217008 184152
rect 216862 181384 216918 181393
rect 216862 181319 216918 181328
rect 216770 81968 216826 81977
rect 216770 81903 216826 81912
rect 216680 66156 216732 66162
rect 216680 66098 216732 66104
rect 216876 65793 216904 181319
rect 216968 69601 216996 184146
rect 217060 73001 217088 185807
rect 217152 78810 217180 192578
rect 217322 184376 217378 184385
rect 217322 184311 217378 184320
rect 217230 183424 217286 183433
rect 217230 183359 217286 183368
rect 217140 78804 217192 78810
rect 217140 78746 217192 78752
rect 217244 77081 217272 183359
rect 217336 78713 217364 184311
rect 217416 181552 217468 181558
rect 217416 181494 217468 181500
rect 217428 80753 217456 181494
rect 217508 151224 217560 151230
rect 217508 151166 217560 151172
rect 217414 80744 217470 80753
rect 217414 80679 217470 80688
rect 217322 78704 217378 78713
rect 217322 78639 217378 78648
rect 217230 77072 217286 77081
rect 217230 77007 217286 77016
rect 217046 72992 217102 73001
rect 217046 72927 217102 72936
rect 216954 69592 217010 69601
rect 216954 69527 217010 69536
rect 217520 67590 217548 151166
rect 218072 72350 218100 195463
rect 218518 188320 218574 188329
rect 218518 188255 218574 188264
rect 218428 185700 218480 185706
rect 218428 185642 218480 185648
rect 218150 183288 218206 183297
rect 218150 183223 218206 183232
rect 218060 72344 218112 72350
rect 218060 72286 218112 72292
rect 217508 67584 217560 67590
rect 217508 67526 217560 67532
rect 218164 66065 218192 183223
rect 218242 183152 218298 183161
rect 218242 183087 218298 183096
rect 218256 182617 218284 183087
rect 218242 182608 218298 182617
rect 218298 182566 218376 182594
rect 218242 182543 218298 182552
rect 218244 182504 218296 182510
rect 218244 182446 218296 182452
rect 218256 70961 218284 182446
rect 218242 70952 218298 70961
rect 218242 70887 218298 70896
rect 218348 69562 218376 182566
rect 218440 182510 218468 185642
rect 218428 182504 218480 182510
rect 218428 182446 218480 182452
rect 218532 182322 218560 188255
rect 218440 182294 218560 182322
rect 218440 76974 218468 182294
rect 218520 181620 218572 181626
rect 218520 181562 218572 181568
rect 218428 76968 218480 76974
rect 218532 76945 218560 181562
rect 218428 76910 218480 76916
rect 218518 76936 218574 76945
rect 218518 76871 218574 76880
rect 218336 69556 218388 69562
rect 218336 69498 218388 69504
rect 218150 66056 218206 66065
rect 218150 65991 218206 66000
rect 216862 65784 216918 65793
rect 216862 65719 216918 65728
rect 216680 65680 216732 65686
rect 216680 65622 216732 65628
rect 215668 46912 215720 46918
rect 215668 46854 215720 46860
rect 216036 46912 216088 46918
rect 216036 46854 216088 46860
rect 215680 46306 215708 46854
rect 215668 46300 215720 46306
rect 215668 46242 215720 46248
rect 216692 16574 216720 65622
rect 219452 62898 219480 198018
rect 219544 63306 219572 198086
rect 220096 195673 220124 699654
rect 220728 198144 220780 198150
rect 220728 198086 220780 198092
rect 220740 197402 220768 198086
rect 220728 197396 220780 197402
rect 220728 197338 220780 197344
rect 220082 195664 220138 195673
rect 220082 195599 220138 195608
rect 224236 192817 224264 699654
rect 230584 683114 230612 703520
rect 230492 683086 230612 683114
rect 230492 271182 230520 683086
rect 230480 271176 230532 271182
rect 230480 271118 230532 271124
rect 224222 192808 224278 192817
rect 224222 192743 224278 192752
rect 219624 183116 219676 183122
rect 219624 183058 219676 183064
rect 219532 63300 219584 63306
rect 219532 63242 219584 63248
rect 219440 62892 219492 62898
rect 219440 62834 219492 62840
rect 219636 52426 219664 183058
rect 219808 183048 219860 183054
rect 219808 182990 219860 182996
rect 219716 180124 219768 180130
rect 219716 180066 219768 180072
rect 219728 60722 219756 180066
rect 219820 66230 219848 182990
rect 233252 181762 233280 703582
rect 234264 703474 234292 703582
rect 234406 703520 234518 704960
rect 237392 703582 238156 703610
rect 234448 703474 234476 703520
rect 234264 703446 234476 703474
rect 237392 194041 237420 703582
rect 238128 703474 238156 703582
rect 238270 703520 238382 704960
rect 241532 703582 242020 703610
rect 238312 703474 238340 703520
rect 238128 703446 238340 703474
rect 237378 194032 237434 194041
rect 237378 193967 237434 193976
rect 241532 188426 241560 703582
rect 241992 703474 242020 703582
rect 242134 703520 242246 704960
rect 245354 703520 245466 704960
rect 249218 703520 249330 704960
rect 253082 703520 253194 704960
rect 256946 703520 257058 704960
rect 260810 703520 260922 704960
rect 264674 703520 264786 704960
rect 268538 703520 268650 704960
rect 272402 703520 272514 704960
rect 276266 703520 276378 704960
rect 280130 703520 280242 704960
rect 283994 703520 284106 704960
rect 287858 703520 287970 704960
rect 291722 703520 291834 704960
rect 295586 703520 295698 704960
rect 299450 703520 299562 704960
rect 302252 703582 302556 703610
rect 242176 703474 242204 703520
rect 241992 703446 242204 703474
rect 245396 699718 245424 703520
rect 249260 702434 249288 703520
rect 253124 702434 253152 703520
rect 256988 702434 257016 703520
rect 248432 702406 249288 702434
rect 252572 702406 253152 702434
rect 256712 702406 257016 702434
rect 242164 699712 242216 699718
rect 242164 699654 242216 699660
rect 245384 699712 245436 699718
rect 245384 699654 245436 699660
rect 242176 189009 242204 699654
rect 242162 189000 242218 189009
rect 242162 188935 242218 188944
rect 241520 188420 241572 188426
rect 241520 188362 241572 188368
rect 248432 185774 248460 702406
rect 252572 200870 252600 702406
rect 252560 200864 252612 200870
rect 252560 200806 252612 200812
rect 256712 191758 256740 702406
rect 256700 191752 256752 191758
rect 256700 191694 256752 191700
rect 260852 189922 260880 703520
rect 264716 702434 264744 703520
rect 268580 702434 268608 703520
rect 263612 702406 264744 702434
rect 267752 702406 268608 702434
rect 263612 268433 263640 702406
rect 263598 268424 263654 268433
rect 263598 268359 263654 268368
rect 267752 263158 267780 702406
rect 272444 699718 272472 703520
rect 276308 702434 276336 703520
rect 276032 702406 276336 702434
rect 269764 699712 269816 699718
rect 269764 699654 269816 699660
rect 272432 699712 272484 699718
rect 272432 699654 272484 699660
rect 267740 263152 267792 263158
rect 267740 263094 267792 263100
rect 260840 189916 260892 189922
rect 260840 189858 260892 189864
rect 269776 188766 269804 699654
rect 276032 263090 276060 702406
rect 280172 699718 280200 703520
rect 284036 702434 284064 703520
rect 282932 702406 284064 702434
rect 278044 699712 278096 699718
rect 278044 699654 278096 699660
rect 280160 699712 280212 699718
rect 280160 699654 280212 699660
rect 276020 263084 276072 263090
rect 276020 263026 276072 263032
rect 269764 188760 269816 188766
rect 269764 188702 269816 188708
rect 278056 187066 278084 699654
rect 278044 187060 278096 187066
rect 278044 187002 278096 187008
rect 282932 186289 282960 702406
rect 287900 700466 287928 703520
rect 291764 702434 291792 703520
rect 291212 702406 291792 702434
rect 287888 700460 287940 700466
rect 287888 700402 287940 700408
rect 291212 199306 291240 702406
rect 299492 262954 299520 703520
rect 299480 262948 299532 262954
rect 299480 262890 299532 262896
rect 302252 199646 302280 703582
rect 302528 703474 302556 703582
rect 302670 703520 302782 704960
rect 306534 703520 306646 704960
rect 310398 703520 310510 704960
rect 313292 703582 314148 703610
rect 302712 703474 302740 703520
rect 302528 703446 302740 703474
rect 306576 683114 306604 703520
rect 310440 703050 310468 703520
rect 309140 703044 309192 703050
rect 309140 702986 309192 702992
rect 310428 703044 310480 703050
rect 310428 702986 310480 702992
rect 306392 683086 306604 683114
rect 302240 199640 302292 199646
rect 302240 199582 302292 199588
rect 291200 199300 291252 199306
rect 291200 199242 291252 199248
rect 282918 186280 282974 186289
rect 282918 186215 282974 186224
rect 248420 185768 248472 185774
rect 248420 185710 248472 185716
rect 306392 185706 306420 683086
rect 306380 185700 306432 185706
rect 306380 185642 306432 185648
rect 309152 182753 309180 702986
rect 313292 183054 313320 703582
rect 314120 703474 314148 703582
rect 314262 703520 314374 704960
rect 318126 703520 318238 704960
rect 321572 703582 321876 703610
rect 314304 703474 314332 703520
rect 314120 703446 314332 703474
rect 313280 183048 313332 183054
rect 313280 182990 313332 182996
rect 309138 182744 309194 182753
rect 309138 182679 309194 182688
rect 233240 181756 233292 181762
rect 233240 181698 233292 181704
rect 321572 179110 321600 703582
rect 321848 703474 321876 703582
rect 321990 703520 322102 704960
rect 325854 703520 325966 704960
rect 329718 703520 329830 704960
rect 332612 703582 333468 703610
rect 322032 703474 322060 703520
rect 321848 703446 322060 703474
rect 325896 699718 325924 703520
rect 329760 703050 329788 703520
rect 328460 703044 328512 703050
rect 328460 702986 328512 702992
rect 329748 703044 329800 703050
rect 329748 702986 329800 702992
rect 323584 699712 323636 699718
rect 323584 699654 323636 699660
rect 325884 699712 325936 699718
rect 325884 699654 325936 699660
rect 323596 195430 323624 699654
rect 323584 195424 323636 195430
rect 323584 195366 323636 195372
rect 328472 193662 328500 702986
rect 328460 193656 328512 193662
rect 328460 193598 328512 193604
rect 332612 192710 332640 703582
rect 333440 703474 333468 703582
rect 333582 703520 333694 704960
rect 337446 703520 337558 704960
rect 340892 703582 341196 703610
rect 333624 703474 333652 703520
rect 333440 703446 333652 703474
rect 340892 194313 340920 703582
rect 341168 703474 341196 703582
rect 341310 703520 341422 704960
rect 345174 703520 345286 704960
rect 349038 703520 349150 704960
rect 351932 703582 352788 703610
rect 341352 703474 341380 703520
rect 341168 703446 341380 703474
rect 349080 703050 349108 703520
rect 347780 703044 347832 703050
rect 347780 702986 347832 702992
rect 349068 703044 349120 703050
rect 349068 702986 349120 702992
rect 347792 263022 347820 702986
rect 347780 263016 347832 263022
rect 347780 262958 347832 262964
rect 340878 194304 340934 194313
rect 340878 194239 340934 194248
rect 332600 192704 332652 192710
rect 332600 192646 332652 192652
rect 321560 179104 321612 179110
rect 321560 179046 321612 179052
rect 351932 175953 351960 703582
rect 352760 703474 352788 703582
rect 352902 703520 353014 704960
rect 356122 703520 356234 704960
rect 359986 703520 360098 704960
rect 363850 703520 363962 704960
rect 367714 703520 367826 704960
rect 371578 703520 371690 704960
rect 375442 703520 375554 704960
rect 379306 703520 379418 704960
rect 383170 703520 383282 704960
rect 387034 703520 387146 704960
rect 390898 703520 391010 704960
rect 394762 703520 394874 704960
rect 398626 703520 398738 704960
rect 402490 703520 402602 704960
rect 406354 703520 406466 704960
rect 410218 703520 410330 704960
rect 412652 703582 413324 703610
rect 352944 703474 352972 703520
rect 352760 703446 352972 703474
rect 356164 683114 356192 703520
rect 360028 703050 360056 703520
rect 358820 703044 358872 703050
rect 358820 702986 358872 702992
rect 360016 703044 360068 703050
rect 360016 702986 360068 702992
rect 356072 683086 356192 683114
rect 356072 181694 356100 683086
rect 356060 181688 356112 181694
rect 356060 181630 356112 181636
rect 358832 177818 358860 702986
rect 363892 702434 363920 703520
rect 367756 702434 367784 703520
rect 371620 702434 371648 703520
rect 362972 702406 363920 702434
rect 367112 702406 367784 702434
rect 371252 702406 371648 702434
rect 362972 180470 363000 702406
rect 362960 180464 363012 180470
rect 362960 180406 363012 180412
rect 358820 177812 358872 177818
rect 358820 177754 358872 177760
rect 367112 176089 367140 702406
rect 371252 189961 371280 702406
rect 375484 699718 375512 703520
rect 379348 703050 379376 703520
rect 378140 703044 378192 703050
rect 378140 702986 378192 702992
rect 379336 703044 379388 703050
rect 379336 702986 379388 702992
rect 374644 699712 374696 699718
rect 374644 699654 374696 699660
rect 375472 699712 375524 699718
rect 375472 699654 375524 699660
rect 374656 201113 374684 699654
rect 374642 201104 374698 201113
rect 374642 201039 374698 201048
rect 371238 189952 371294 189961
rect 371238 189887 371294 189896
rect 378152 188465 378180 702986
rect 383212 702434 383240 703520
rect 387076 702434 387104 703520
rect 382292 702406 383240 702434
rect 386432 702406 387104 702434
rect 378138 188456 378194 188465
rect 378138 188391 378194 188400
rect 382292 176225 382320 702406
rect 386432 195809 386460 702406
rect 394804 700398 394832 703520
rect 394792 700392 394844 700398
rect 394792 700334 394844 700340
rect 398668 699718 398696 703520
rect 402532 699718 402560 703520
rect 406396 702434 406424 703520
rect 410260 702434 410288 703520
rect 405752 702406 406424 702434
rect 409892 702406 410288 702434
rect 395344 699712 395396 699718
rect 395344 699654 395396 699660
rect 398656 699712 398708 699718
rect 398656 699654 398708 699660
rect 400864 699712 400916 699718
rect 400864 699654 400916 699660
rect 402520 699712 402572 699718
rect 402520 699654 402572 699660
rect 386418 195800 386474 195809
rect 386418 195735 386474 195744
rect 395356 176526 395384 699654
rect 400876 264246 400904 699654
rect 400864 264240 400916 264246
rect 400864 264182 400916 264188
rect 405752 179178 405780 702406
rect 409892 183569 409920 702406
rect 412652 199510 412680 703582
rect 413296 703474 413324 703582
rect 413438 703520 413550 704960
rect 416792 703582 417188 703610
rect 413480 703474 413508 703520
rect 413296 703446 413508 703474
rect 412640 199504 412692 199510
rect 412640 199446 412692 199452
rect 416792 191593 416820 703582
rect 417160 703474 417188 703582
rect 417302 703520 417414 704960
rect 421166 703520 421278 704960
rect 425030 703520 425142 704960
rect 427832 703582 428780 703610
rect 417344 703474 417372 703520
rect 417160 703446 417372 703474
rect 421208 702434 421236 703520
rect 420932 702406 421236 702434
rect 420932 196897 420960 702406
rect 420918 196888 420974 196897
rect 420918 196823 420974 196832
rect 425072 194449 425100 703520
rect 427832 199578 427860 703582
rect 428752 703474 428780 703582
rect 428894 703520 429006 704960
rect 431972 703582 432644 703610
rect 428936 703474 428964 703520
rect 428752 703446 428964 703474
rect 427820 199572 427872 199578
rect 427820 199514 427872 199520
rect 431972 199442 432000 703582
rect 432616 703474 432644 703582
rect 432758 703520 432870 704960
rect 436112 703582 436508 703610
rect 432800 703474 432828 703520
rect 432616 703446 432828 703474
rect 431960 199436 432012 199442
rect 431960 199378 432012 199384
rect 425058 194440 425114 194449
rect 425058 194375 425114 194384
rect 416778 191584 416834 191593
rect 416778 191519 416834 191528
rect 436112 184278 436140 703582
rect 436480 703474 436508 703582
rect 436622 703520 436734 704960
rect 440486 703520 440598 704960
rect 444350 703520 444462 704960
rect 448214 703520 448326 704960
rect 452078 703520 452190 704960
rect 455432 703582 455828 703610
rect 436664 703474 436692 703520
rect 436480 703446 436692 703474
rect 440528 702434 440556 703520
rect 440252 702406 440556 702434
rect 440252 191457 440280 702406
rect 440238 191448 440294 191457
rect 440238 191383 440294 191392
rect 444392 184521 444420 703520
rect 448256 699718 448284 703520
rect 452120 699718 452148 703520
rect 445024 699712 445076 699718
rect 445024 699654 445076 699660
rect 448244 699712 448296 699718
rect 448244 699654 448296 699660
rect 449164 699712 449216 699718
rect 449164 699654 449216 699660
rect 452108 699712 452160 699718
rect 452108 699654 452160 699660
rect 445036 197169 445064 699654
rect 445022 197160 445078 197169
rect 445022 197095 445078 197104
rect 449176 188834 449204 699654
rect 449164 188828 449216 188834
rect 449164 188770 449216 188776
rect 444378 184512 444434 184521
rect 444378 184447 444434 184456
rect 436100 184272 436152 184278
rect 436100 184214 436152 184220
rect 409878 183560 409934 183569
rect 409878 183495 409934 183504
rect 455432 180538 455460 703582
rect 455800 703474 455828 703582
rect 455942 703520 456054 704960
rect 459806 703520 459918 704960
rect 463670 703520 463782 704960
rect 466472 703582 467420 703610
rect 455984 703474 456012 703520
rect 455800 703446 456012 703474
rect 459848 702434 459876 703520
rect 459572 702406 459876 702434
rect 459572 182073 459600 702406
rect 463712 183433 463740 703520
rect 466472 201793 466500 703582
rect 467392 703474 467420 703582
rect 467534 703520 467646 704960
rect 470754 703520 470866 704960
rect 474618 703520 474730 704960
rect 478482 703520 478594 704960
rect 482346 703520 482458 704960
rect 486210 703520 486322 704960
rect 490074 703520 490186 704960
rect 493938 703520 494050 704960
rect 497802 703520 497914 704960
rect 501666 703520 501778 704960
rect 505530 703520 505642 704960
rect 509394 703520 509506 704960
rect 513258 703520 513370 704960
rect 517122 703520 517234 704960
rect 520986 703520 521098 704960
rect 524850 703520 524962 704960
rect 527192 703582 527956 703610
rect 467576 703474 467604 703520
rect 467392 703446 467604 703474
rect 470796 683114 470824 703520
rect 474660 699718 474688 703520
rect 478524 702434 478552 703520
rect 482388 702434 482416 703520
rect 486252 702434 486280 703520
rect 477512 702406 478552 702434
rect 481652 702406 482416 702434
rect 485792 702406 486280 702434
rect 472624 699712 472676 699718
rect 472624 699654 472676 699660
rect 474648 699712 474700 699718
rect 474648 699654 474700 699660
rect 470612 683086 470824 683114
rect 470612 263566 470640 683086
rect 472636 268394 472664 699654
rect 472624 268388 472676 268394
rect 472624 268330 472676 268336
rect 470600 263560 470652 263566
rect 470600 263502 470652 263508
rect 477512 262886 477540 702406
rect 477500 262880 477552 262886
rect 477500 262822 477552 262828
rect 466458 201784 466514 201793
rect 466458 201719 466514 201728
rect 463698 183424 463754 183433
rect 463698 183359 463754 183368
rect 459558 182064 459614 182073
rect 459558 181999 459614 182008
rect 455420 180532 455472 180538
rect 455420 180474 455472 180480
rect 481652 180305 481680 702406
rect 485792 195945 485820 702406
rect 490116 683114 490144 703520
rect 493980 697610 494008 703520
rect 497844 699718 497872 703520
rect 501708 699718 501736 703520
rect 505572 699718 505600 703520
rect 494704 699712 494756 699718
rect 494704 699654 494756 699660
rect 497832 699712 497884 699718
rect 497832 699654 497884 699660
rect 498844 699712 498896 699718
rect 498844 699654 498896 699660
rect 501696 699712 501748 699718
rect 501696 699654 501748 699660
rect 502984 699712 503036 699718
rect 502984 699654 503036 699660
rect 505560 699712 505612 699718
rect 505560 699654 505612 699660
rect 492680 697604 492732 697610
rect 492680 697546 492732 697552
rect 493968 697604 494020 697610
rect 493968 697546 494020 697552
rect 489932 683086 490144 683114
rect 485778 195936 485834 195945
rect 485778 195871 485834 195880
rect 489932 183297 489960 683086
rect 492692 265674 492720 697546
rect 492680 265668 492732 265674
rect 492680 265610 492732 265616
rect 489918 183288 489974 183297
rect 489918 183223 489974 183232
rect 494716 180441 494744 699654
rect 498856 278050 498884 699654
rect 498844 278044 498896 278050
rect 498844 277986 498896 277992
rect 498844 260908 498896 260914
rect 498844 260850 498896 260856
rect 498856 238746 498884 260850
rect 498844 238740 498896 238746
rect 498844 238682 498896 238688
rect 502996 194002 503024 699654
rect 509436 683114 509464 703520
rect 513300 697610 513328 703520
rect 517164 702434 517192 703520
rect 521028 702434 521056 703520
rect 524892 702434 524920 703520
rect 516152 702406 517192 702434
rect 520292 702406 521056 702434
rect 524432 702406 524920 702434
rect 512000 697604 512052 697610
rect 512000 697546 512052 697552
rect 513288 697604 513340 697610
rect 513288 697546 513340 697552
rect 509252 683086 509464 683114
rect 509252 200977 509280 683086
rect 509238 200968 509294 200977
rect 509238 200903 509294 200912
rect 502984 193996 503036 194002
rect 502984 193938 503036 193944
rect 512012 186182 512040 697546
rect 516152 191321 516180 702406
rect 520292 262721 520320 702406
rect 524432 276690 524460 702406
rect 524420 276684 524472 276690
rect 524420 276626 524472 276632
rect 520278 262712 520334 262721
rect 520278 262647 520334 262656
rect 516138 191312 516194 191321
rect 516138 191247 516194 191256
rect 527192 188358 527220 703582
rect 527928 703474 527956 703582
rect 528070 703520 528182 704960
rect 531934 703520 532046 704960
rect 535472 703582 535684 703610
rect 528112 703474 528140 703520
rect 527928 703446 528140 703474
rect 535472 269793 535500 703582
rect 535656 703474 535684 703582
rect 535798 703520 535910 704960
rect 539662 703520 539774 704960
rect 542372 703582 543412 703610
rect 535840 703474 535868 703520
rect 535656 703446 535868 703474
rect 539704 683114 539732 703520
rect 539612 683086 539732 683114
rect 535458 269784 535514 269793
rect 535458 269719 535514 269728
rect 527180 188352 527232 188358
rect 527180 188294 527232 188300
rect 512000 186176 512052 186182
rect 512000 186118 512052 186124
rect 539612 181393 539640 683086
rect 542372 194585 542400 703582
rect 543384 703474 543412 703582
rect 543526 703520 543638 704960
rect 546512 703582 547276 703610
rect 543568 703474 543596 703520
rect 543384 703446 543596 703474
rect 544384 694204 544436 694210
rect 544384 694146 544436 694152
rect 542358 194576 542414 194585
rect 542358 194511 542414 194520
rect 539598 181384 539654 181393
rect 539598 181319 539654 181328
rect 494702 180432 494758 180441
rect 494702 180367 494758 180376
rect 481638 180296 481694 180305
rect 481638 180231 481694 180240
rect 405740 179172 405792 179178
rect 405740 179114 405792 179120
rect 395344 176520 395396 176526
rect 395344 176462 395396 176468
rect 544396 176361 544424 694146
rect 544476 568608 544528 568614
rect 544476 568550 544528 568556
rect 544488 177993 544516 568550
rect 546512 188329 546540 703582
rect 547248 703474 547276 703582
rect 547390 703520 547502 704960
rect 551254 703520 551366 704960
rect 555118 703520 555230 704960
rect 558982 703520 559094 704960
rect 561692 703582 562732 703610
rect 547432 703474 547460 703520
rect 547248 703446 547460 703474
rect 548616 700392 548668 700398
rect 548616 700334 548668 700340
rect 548524 685908 548576 685914
rect 548524 685850 548576 685856
rect 546498 188320 546554 188329
rect 546498 188255 546554 188264
rect 544474 177984 544530 177993
rect 544474 177919 544530 177928
rect 548536 176633 548564 685850
rect 548628 199617 548656 700334
rect 551296 700330 551324 703520
rect 551284 700324 551336 700330
rect 551284 700266 551336 700272
rect 555160 699718 555188 703520
rect 556804 700324 556856 700330
rect 556804 700266 556856 700272
rect 552664 699712 552716 699718
rect 552664 699654 552716 699660
rect 555148 699712 555200 699718
rect 555148 699654 555200 699660
rect 548614 199608 548670 199617
rect 548614 199543 548670 199552
rect 552676 184249 552704 699654
rect 552756 629332 552808 629338
rect 552756 629274 552808 629280
rect 552662 184240 552718 184249
rect 552662 184175 552718 184184
rect 552768 181490 552796 629274
rect 554044 543788 554096 543794
rect 554044 543730 554096 543736
rect 552848 459604 552900 459610
rect 552848 459546 552900 459552
rect 552756 181484 552808 181490
rect 552756 181426 552808 181432
rect 552860 176662 552888 459546
rect 554056 177954 554084 543730
rect 555424 371272 555476 371278
rect 555424 371214 555476 371220
rect 555436 178022 555464 371214
rect 555516 282940 555568 282946
rect 555516 282882 555568 282888
rect 555424 178016 555476 178022
rect 555424 177958 555476 177964
rect 554044 177948 554096 177954
rect 554044 177890 554096 177896
rect 552848 176656 552900 176662
rect 548522 176624 548578 176633
rect 552848 176598 552900 176604
rect 555528 176594 555556 282882
rect 556816 180742 556844 700266
rect 559024 683114 559052 703520
rect 558932 683086 559052 683114
rect 556896 669384 556948 669390
rect 556896 669326 556948 669332
rect 556804 180736 556856 180742
rect 556804 180678 556856 180684
rect 556908 178673 556936 669326
rect 558184 507884 558236 507890
rect 558184 507826 558236 507832
rect 558196 179246 558224 507826
rect 558276 495508 558328 495514
rect 558276 495450 558328 495456
rect 558184 179240 558236 179246
rect 558184 179182 558236 179188
rect 556894 178664 556950 178673
rect 556894 178599 556950 178608
rect 548522 176559 548578 176568
rect 555516 176588 555568 176594
rect 555516 176530 555568 176536
rect 558288 176497 558316 495450
rect 558368 455456 558420 455462
rect 558368 455398 558420 455404
rect 558380 180606 558408 455398
rect 558460 310548 558512 310554
rect 558460 310490 558512 310496
rect 558472 186250 558500 310490
rect 558552 289876 558604 289882
rect 558552 289818 558604 289824
rect 558460 186244 558512 186250
rect 558460 186186 558512 186192
rect 558564 180674 558592 289818
rect 558932 195129 558960 683086
rect 560944 527196 560996 527202
rect 560944 527138 560996 527144
rect 558918 195120 558974 195129
rect 558918 195055 558974 195064
rect 558552 180668 558604 180674
rect 558552 180610 558604 180616
rect 558368 180600 558420 180606
rect 558368 180542 558420 180548
rect 560956 178702 560984 527138
rect 561036 474768 561088 474774
rect 561036 474710 561088 474716
rect 561048 184385 561076 474710
rect 561128 472048 561180 472054
rect 561128 471990 561180 471996
rect 561140 192642 561168 471990
rect 561220 443012 561272 443018
rect 561220 442954 561272 442960
rect 561128 192636 561180 192642
rect 561128 192578 561180 192584
rect 561034 184376 561090 184385
rect 561034 184311 561090 184320
rect 561232 182170 561260 442954
rect 561312 278792 561364 278798
rect 561312 278734 561364 278740
rect 561324 198014 561352 278734
rect 561692 200841 561720 703582
rect 562704 703474 562732 703582
rect 562846 703520 562958 704960
rect 566710 703520 566822 704960
rect 570574 703520 570686 704960
rect 574438 703520 574550 704960
rect 578302 703520 578414 704960
rect 581012 703582 582052 703610
rect 562888 703474 562916 703520
rect 562704 703446 562916 703474
rect 570616 700398 570644 703520
rect 570604 700392 570656 700398
rect 570604 700334 570656 700340
rect 574480 700330 574508 703520
rect 576124 702500 576176 702506
rect 576124 702442 576176 702448
rect 574468 700324 574520 700330
rect 574468 700266 574520 700272
rect 570604 698352 570656 698358
rect 570604 698294 570656 698300
rect 566464 644496 566516 644502
rect 566464 644438 566516 644444
rect 565084 608660 565136 608666
rect 565084 608602 565136 608608
rect 562324 523048 562376 523054
rect 562324 522990 562376 522996
rect 561678 200832 561734 200841
rect 561678 200767 561734 200776
rect 562336 200734 562364 522990
rect 563704 478916 563756 478922
rect 563704 478858 563756 478864
rect 562416 463752 562468 463758
rect 562416 463694 562468 463700
rect 562324 200728 562376 200734
rect 562324 200670 562376 200676
rect 561312 198008 561364 198014
rect 561312 197950 561364 197956
rect 561220 182164 561272 182170
rect 561220 182106 561272 182112
rect 562428 181626 562456 463694
rect 563716 196654 563744 478858
rect 563796 467900 563848 467906
rect 563796 467842 563848 467848
rect 563704 196648 563756 196654
rect 563704 196590 563756 196596
rect 563808 188902 563836 467842
rect 563888 426488 563940 426494
rect 563888 426430 563940 426436
rect 563796 188896 563848 188902
rect 563796 188838 563848 188844
rect 563900 184210 563928 426430
rect 563980 342304 564032 342310
rect 563980 342246 564032 342252
rect 563888 184204 563940 184210
rect 563888 184146 563940 184152
rect 562416 181620 562468 181626
rect 562416 181562 562468 181568
rect 563992 180810 564020 342246
rect 564072 306400 564124 306406
rect 564072 306342 564124 306348
rect 564084 181558 564112 306342
rect 565096 183025 565124 608602
rect 565176 403028 565228 403034
rect 565176 402970 565228 402976
rect 565082 183016 565138 183025
rect 565082 182951 565138 182960
rect 564072 181552 564124 181558
rect 564072 181494 564124 181500
rect 563980 180804 564032 180810
rect 563980 180746 564032 180752
rect 565188 180577 565216 402970
rect 566476 187377 566504 644438
rect 567844 633480 567896 633486
rect 567844 633422 567896 633428
rect 566648 572756 566700 572762
rect 566648 572698 566700 572704
rect 566556 512032 566608 512038
rect 566556 511974 566608 511980
rect 566568 189825 566596 511974
rect 566554 189816 566610 189825
rect 566554 189751 566610 189760
rect 566660 187513 566688 572698
rect 566740 358828 566792 358834
rect 566740 358770 566792 358776
rect 566646 187504 566702 187513
rect 566646 187439 566702 187448
rect 566462 187368 566518 187377
rect 566462 187303 566518 187312
rect 566752 185638 566780 358770
rect 566832 274712 566884 274718
rect 566832 274654 566884 274660
rect 566740 185632 566792 185638
rect 566740 185574 566792 185580
rect 566844 182986 566872 274654
rect 567856 191185 567884 633422
rect 567936 596216 567988 596222
rect 567936 596158 567988 596164
rect 567842 191176 567898 191185
rect 567842 191111 567898 191120
rect 567948 185881 567976 596158
rect 569224 487212 569276 487218
rect 569224 487154 569276 487160
rect 568028 430636 568080 430642
rect 568028 430578 568080 430584
rect 568040 188970 568068 430578
rect 568028 188964 568080 188970
rect 568028 188906 568080 188912
rect 569236 187678 569264 487154
rect 569316 346452 569368 346458
rect 569316 346394 569368 346400
rect 569224 187672 569276 187678
rect 569224 187614 569276 187620
rect 569328 186969 569356 346394
rect 569408 302252 569460 302258
rect 569408 302194 569460 302200
rect 569314 186960 569370 186969
rect 569314 186895 569370 186904
rect 569420 186318 569448 302194
rect 570616 189038 570644 698294
rect 574744 583772 574796 583778
rect 574744 583714 574796 583720
rect 571984 564460 572036 564466
rect 571984 564402 572036 564408
rect 570696 539640 570748 539646
rect 570696 539582 570748 539588
rect 570604 189032 570656 189038
rect 570604 188974 570656 188980
rect 569408 186312 569460 186318
rect 569408 186254 569460 186260
rect 567934 185872 567990 185881
rect 567934 185807 567990 185816
rect 566832 182980 566884 182986
rect 566832 182922 566884 182928
rect 565174 180568 565230 180577
rect 565174 180503 565230 180512
rect 570708 178945 570736 539582
rect 570788 434784 570840 434790
rect 570788 434726 570840 434732
rect 570800 185745 570828 434726
rect 571996 195401 572024 564402
rect 573364 516180 573416 516186
rect 573364 516122 573416 516128
rect 572076 447160 572128 447166
rect 572076 447102 572128 447108
rect 571982 195392 572038 195401
rect 571982 195327 572038 195336
rect 572088 186998 572116 447102
rect 572168 390584 572220 390590
rect 572168 390526 572220 390532
rect 572180 187241 572208 390526
rect 572260 331288 572312 331294
rect 572260 331230 572312 331236
rect 572272 189854 572300 331230
rect 572352 285728 572404 285734
rect 572352 285670 572404 285676
rect 572260 189848 572312 189854
rect 572260 189790 572312 189796
rect 572166 187232 572222 187241
rect 572166 187167 572222 187176
rect 572076 186992 572128 186998
rect 572076 186934 572128 186940
rect 570786 185736 570842 185745
rect 570786 185671 570842 185680
rect 572364 184822 572392 285670
rect 572352 184816 572404 184822
rect 572352 184758 572404 184764
rect 570694 178936 570750 178945
rect 570694 178871 570750 178880
rect 573376 178809 573404 516122
rect 574756 195362 574784 583714
rect 574836 520328 574888 520334
rect 574836 520270 574888 520276
rect 574744 195356 574796 195362
rect 574744 195298 574796 195304
rect 574848 192681 574876 520270
rect 574928 423700 574980 423706
rect 574928 423642 574980 423648
rect 574834 192672 574890 192681
rect 574834 192607 574890 192616
rect 574940 190369 574968 423642
rect 575112 411324 575164 411330
rect 575112 411266 575164 411272
rect 575020 314696 575072 314702
rect 575020 314638 575072 314644
rect 574926 190360 574982 190369
rect 574926 190295 574982 190304
rect 575032 187105 575060 314638
rect 575124 189689 575152 411266
rect 576136 196761 576164 702442
rect 578344 683114 578372 703520
rect 580170 702536 580226 702545
rect 580170 702471 580172 702480
rect 580224 702471 580226 702480
rect 580172 702442 580224 702448
rect 580170 698456 580226 698465
rect 580170 698391 580226 698400
rect 580184 698358 580212 698391
rect 580172 698352 580224 698358
rect 580172 698294 580224 698300
rect 580170 694376 580226 694385
rect 580170 694311 580226 694320
rect 580184 694210 580212 694311
rect 580172 694204 580224 694210
rect 580172 694146 580224 694152
rect 579802 686216 579858 686225
rect 579802 686151 579858 686160
rect 579816 685914 579844 686151
rect 579804 685908 579856 685914
rect 579804 685850 579856 685856
rect 578252 683086 578372 683114
rect 576216 677612 576268 677618
rect 576216 677554 576268 677560
rect 576122 196752 576178 196761
rect 576122 196687 576178 196696
rect 576228 191049 576256 677554
rect 577504 625456 577556 625462
rect 577504 625398 577556 625404
rect 576308 499588 576360 499594
rect 576308 499530 576360 499536
rect 576320 196625 576348 499530
rect 576400 394732 576452 394738
rect 576400 394674 576452 394680
rect 576306 196616 576362 196625
rect 576306 196551 576362 196560
rect 576412 193118 576440 394674
rect 577516 195265 577544 625398
rect 577596 338156 577648 338162
rect 577596 338098 577648 338104
rect 577502 195256 577558 195265
rect 577502 195191 577558 195200
rect 576400 193112 576452 193118
rect 576400 193054 576452 193060
rect 577608 193050 577636 338098
rect 577688 318844 577740 318850
rect 577688 318786 577740 318792
rect 577596 193044 577648 193050
rect 577596 192986 577648 192992
rect 576214 191040 576270 191049
rect 576214 190975 576270 190984
rect 577700 190398 577728 318786
rect 577872 270564 577924 270570
rect 577872 270506 577924 270512
rect 577780 262268 577832 262274
rect 577780 262210 577832 262216
rect 577688 190392 577740 190398
rect 577688 190334 577740 190340
rect 575110 189680 575166 189689
rect 575110 189615 575166 189624
rect 575018 187096 575074 187105
rect 575018 187031 575074 187040
rect 573362 178800 573418 178809
rect 577792 178770 577820 262210
rect 577884 192506 577912 270506
rect 578252 192545 578280 683086
rect 580170 678056 580226 678065
rect 580170 677991 580226 678000
rect 580184 677618 580212 677991
rect 580172 677612 580224 677618
rect 580172 677554 580224 677560
rect 580170 669896 580226 669905
rect 580170 669831 580226 669840
rect 580184 669390 580212 669831
rect 580172 669384 580224 669390
rect 580172 669326 580224 669332
rect 580170 665816 580226 665825
rect 580170 665751 580226 665760
rect 580184 665242 580212 665751
rect 580172 665236 580224 665242
rect 580172 665178 580224 665184
rect 579986 649496 580042 649505
rect 579986 649431 580042 649440
rect 580000 648650 580028 649431
rect 579988 648644 580040 648650
rect 579988 648586 580040 648592
rect 580170 645416 580226 645425
rect 580170 645351 580226 645360
rect 580184 644502 580212 645351
rect 580172 644496 580224 644502
rect 580172 644438 580224 644444
rect 580170 633856 580226 633865
rect 580170 633791 580226 633800
rect 580184 633486 580212 633791
rect 580172 633480 580224 633486
rect 580172 633422 580224 633428
rect 580170 629776 580226 629785
rect 580170 629711 580226 629720
rect 580184 629338 580212 629711
rect 580172 629332 580224 629338
rect 580172 629274 580224 629280
rect 580538 625696 580594 625705
rect 580538 625631 580594 625640
rect 580552 625462 580580 625631
rect 580540 625456 580592 625462
rect 580540 625398 580592 625404
rect 580170 609376 580226 609385
rect 580170 609311 580226 609320
rect 580184 608666 580212 609311
rect 580172 608660 580224 608666
rect 580172 608602 580224 608608
rect 580354 605296 580410 605305
rect 580354 605231 580410 605240
rect 580170 597136 580226 597145
rect 580170 597071 580226 597080
rect 580184 596222 580212 597071
rect 580172 596216 580224 596222
rect 580172 596158 580224 596164
rect 580170 593056 580226 593065
rect 580170 592991 580226 593000
rect 580184 592074 580212 592991
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 584896 580226 584905
rect 580170 584831 580226 584840
rect 580184 583778 580212 584831
rect 580172 583772 580224 583778
rect 580172 583714 580224 583720
rect 578882 577416 578938 577425
rect 578882 577351 578938 577360
rect 578238 192536 578294 192545
rect 577872 192500 577924 192506
rect 578238 192471 578294 192480
rect 577872 192442 577924 192448
rect 578896 191146 578924 577351
rect 580170 573336 580226 573345
rect 580170 573271 580226 573280
rect 580184 572762 580212 573271
rect 580172 572756 580224 572762
rect 580172 572698 580224 572704
rect 579710 569256 579766 569265
rect 579710 569191 579766 569200
rect 579724 568614 579752 569191
rect 579712 568608 579764 568614
rect 579712 568550 579764 568556
rect 580170 565176 580226 565185
rect 580170 565111 580226 565120
rect 580184 564466 580212 565111
rect 580172 564460 580224 564466
rect 580172 564402 580224 564408
rect 579618 561096 579674 561105
rect 579618 561031 579674 561040
rect 579632 560318 579660 561031
rect 579620 560312 579672 560318
rect 579620 560254 579672 560260
rect 580078 548856 580134 548865
rect 580078 548791 580134 548800
rect 580092 547942 580120 548791
rect 580080 547936 580132 547942
rect 580080 547878 580132 547884
rect 580170 544776 580226 544785
rect 580170 544711 580226 544720
rect 580184 543794 580212 544711
rect 580172 543788 580224 543794
rect 580172 543730 580224 543736
rect 579710 540696 579766 540705
rect 579710 540631 579766 540640
rect 579724 539646 579752 540631
rect 579712 539640 579764 539646
rect 579712 539582 579764 539588
rect 580170 536616 580226 536625
rect 580170 536551 580226 536560
rect 580184 535498 580212 536551
rect 580172 535492 580224 535498
rect 580172 535434 580224 535440
rect 580170 528456 580226 528465
rect 580170 528391 580226 528400
rect 580184 527202 580212 528391
rect 580172 527196 580224 527202
rect 580172 527138 580224 527144
rect 580170 524376 580226 524385
rect 580170 524311 580226 524320
rect 580184 523054 580212 524311
rect 580172 523048 580224 523054
rect 580172 522990 580224 522996
rect 579710 520976 579766 520985
rect 579710 520911 579766 520920
rect 579724 520334 579752 520911
rect 579712 520328 579764 520334
rect 579712 520270 579764 520276
rect 580170 516896 580226 516905
rect 580170 516831 580226 516840
rect 580184 516186 580212 516831
rect 580172 516180 580224 516186
rect 580172 516122 580224 516128
rect 579618 512816 579674 512825
rect 579618 512751 579674 512760
rect 579632 512038 579660 512751
rect 579620 512032 579672 512038
rect 579620 511974 579672 511980
rect 580170 508736 580226 508745
rect 580170 508671 580226 508680
rect 580184 507890 580212 508671
rect 580172 507884 580224 507890
rect 580172 507826 580224 507832
rect 580078 504656 580134 504665
rect 580078 504591 580134 504600
rect 580092 503742 580120 504591
rect 580080 503736 580132 503742
rect 580080 503678 580132 503684
rect 580170 500576 580226 500585
rect 580170 500511 580226 500520
rect 580184 499594 580212 500511
rect 580172 499588 580224 499594
rect 580172 499530 580224 499536
rect 580170 496496 580226 496505
rect 580170 496431 580226 496440
rect 580184 495514 580212 496431
rect 580172 495508 580224 495514
rect 580172 495450 580224 495456
rect 580170 488336 580226 488345
rect 580170 488271 580226 488280
rect 580184 487218 580212 488271
rect 580172 487212 580224 487218
rect 580172 487154 580224 487160
rect 580170 484256 580226 484265
rect 580170 484191 580226 484200
rect 580184 483070 580212 484191
rect 580172 483064 580224 483070
rect 580172 483006 580224 483012
rect 580170 480176 580226 480185
rect 580170 480111 580226 480120
rect 580184 478922 580212 480111
rect 580172 478916 580224 478922
rect 580172 478858 580224 478864
rect 580170 476096 580226 476105
rect 580170 476031 580226 476040
rect 580184 474774 580212 476031
rect 580172 474768 580224 474774
rect 580172 474710 580224 474716
rect 580172 472048 580224 472054
rect 580170 472016 580172 472025
rect 580224 472016 580226 472025
rect 580170 471951 580226 471960
rect 580170 467936 580226 467945
rect 580170 467871 580172 467880
rect 580224 467871 580226 467880
rect 580172 467842 580224 467848
rect 580170 463856 580226 463865
rect 580170 463791 580226 463800
rect 580184 463758 580212 463791
rect 580172 463752 580224 463758
rect 580172 463694 580224 463700
rect 580170 460456 580226 460465
rect 580170 460391 580226 460400
rect 580184 459610 580212 460391
rect 580172 459604 580224 459610
rect 580172 459546 580224 459552
rect 580078 456376 580134 456385
rect 580078 456311 580134 456320
rect 580092 455462 580120 456311
rect 580080 455456 580132 455462
rect 580080 455398 580132 455404
rect 580170 452296 580226 452305
rect 580170 452231 580226 452240
rect 580184 451314 580212 452231
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 579710 448216 579766 448225
rect 579710 448151 579766 448160
rect 579724 447166 579752 448151
rect 579712 447160 579764 447166
rect 579712 447102 579764 447108
rect 580170 444136 580226 444145
rect 580170 444071 580226 444080
rect 580184 443018 580212 444071
rect 580172 443012 580224 443018
rect 580172 442954 580224 442960
rect 580170 435976 580226 435985
rect 580170 435911 580226 435920
rect 580184 434790 580212 435911
rect 580172 434784 580224 434790
rect 580172 434726 580224 434732
rect 580170 431896 580226 431905
rect 580170 431831 580226 431840
rect 580184 430642 580212 431831
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 427816 580226 427825
rect 580170 427751 580226 427760
rect 580184 426494 580212 427751
rect 580172 426488 580224 426494
rect 580172 426430 580224 426436
rect 580170 423736 580226 423745
rect 580170 423671 580172 423680
rect 580224 423671 580226 423680
rect 580172 423642 580224 423648
rect 580170 419656 580226 419665
rect 580170 419591 580226 419600
rect 580184 419558 580212 419591
rect 580172 419552 580224 419558
rect 580172 419494 580224 419500
rect 580170 415576 580226 415585
rect 580170 415511 580226 415520
rect 580184 415478 580212 415511
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 579986 411496 580042 411505
rect 579986 411431 580042 411440
rect 580000 411330 580028 411431
rect 579988 411324 580040 411330
rect 579988 411266 580040 411272
rect 580170 407416 580226 407425
rect 580170 407351 580226 407360
rect 580184 407182 580212 407351
rect 580172 407176 580224 407182
rect 580172 407118 580224 407124
rect 580170 404016 580226 404025
rect 580170 403951 580226 403960
rect 580184 403034 580212 403951
rect 580172 403028 580224 403034
rect 580172 402970 580224 402976
rect 579710 399936 579766 399945
rect 579710 399871 579766 399880
rect 579724 398886 579752 399871
rect 579712 398880 579764 398886
rect 579712 398822 579764 398828
rect 580170 395856 580226 395865
rect 580170 395791 580226 395800
rect 580184 394738 580212 395791
rect 580172 394732 580224 394738
rect 580172 394674 580224 394680
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 580184 390590 580212 391711
rect 580172 390584 580224 390590
rect 580172 390526 580224 390532
rect 580170 387696 580226 387705
rect 580170 387631 580226 387640
rect 580184 386442 580212 387631
rect 580172 386436 580224 386442
rect 580172 386378 580224 386384
rect 578974 383616 579030 383625
rect 578974 383551 579030 383560
rect 578884 191140 578936 191146
rect 578884 191082 578936 191088
rect 578988 179314 579016 383551
rect 580170 375456 580226 375465
rect 580170 375391 580172 375400
rect 580224 375391 580226 375400
rect 580172 375362 580224 375368
rect 579802 371376 579858 371385
rect 579802 371311 579858 371320
rect 579816 371278 579844 371311
rect 579804 371272 579856 371278
rect 579804 371214 579856 371220
rect 580170 367296 580226 367305
rect 580170 367231 580226 367240
rect 580184 367130 580212 367231
rect 580172 367124 580224 367130
rect 580172 367066 580224 367072
rect 580170 359136 580226 359145
rect 580170 359071 580226 359080
rect 580184 358834 580212 359071
rect 580172 358828 580224 358834
rect 580172 358770 580224 358776
rect 580170 355056 580226 355065
rect 580170 354991 580226 355000
rect 580184 354754 580212 354991
rect 580172 354748 580224 354754
rect 580172 354690 580224 354696
rect 580170 350976 580226 350985
rect 580170 350911 580226 350920
rect 580184 350606 580212 350911
rect 580172 350600 580224 350606
rect 580172 350542 580224 350548
rect 580170 346896 580226 346905
rect 580170 346831 580226 346840
rect 580184 346458 580212 346831
rect 580172 346452 580224 346458
rect 580172 346394 580224 346400
rect 579710 343496 579766 343505
rect 579710 343431 579766 343440
rect 579724 342310 579752 343431
rect 579712 342304 579764 342310
rect 579712 342246 579764 342252
rect 579618 339416 579674 339425
rect 579618 339351 579674 339360
rect 579632 338162 579660 339351
rect 579620 338156 579672 338162
rect 579620 338098 579672 338104
rect 579712 331288 579764 331294
rect 579710 331256 579712 331265
rect 579764 331256 579766 331265
rect 579710 331191 579766 331200
rect 579066 323096 579122 323105
rect 579066 323031 579122 323040
rect 579080 189786 579108 323031
rect 579710 319016 579766 319025
rect 579710 318951 579766 318960
rect 579724 318850 579752 318951
rect 579712 318844 579764 318850
rect 579712 318786 579764 318792
rect 579618 314936 579674 314945
rect 579618 314871 579674 314880
rect 579632 314702 579660 314871
rect 579620 314696 579672 314702
rect 579620 314638 579672 314644
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580184 310554 580212 310791
rect 580172 310548 580224 310554
rect 580172 310490 580224 310496
rect 580170 306776 580226 306785
rect 580170 306711 580226 306720
rect 580184 306406 580212 306711
rect 580172 306400 580224 306406
rect 580172 306342 580224 306348
rect 580170 302696 580226 302705
rect 580170 302631 580226 302640
rect 580184 302258 580212 302631
rect 580172 302252 580224 302258
rect 580172 302194 580224 302200
rect 579158 298616 579214 298625
rect 579158 298551 579214 298560
rect 579172 191826 579200 298551
rect 580170 294536 580226 294545
rect 580170 294471 580226 294480
rect 580184 294030 580212 294471
rect 580172 294024 580224 294030
rect 580172 293966 580224 293972
rect 579986 290456 580042 290465
rect 579986 290391 580042 290400
rect 580000 289882 580028 290391
rect 579988 289876 580040 289882
rect 579988 289818 580040 289824
rect 579986 286376 580042 286385
rect 579986 286311 580042 286320
rect 580000 285734 580028 286311
rect 579988 285728 580040 285734
rect 579988 285670 580040 285676
rect 580170 282976 580226 282985
rect 580170 282911 580172 282920
rect 580224 282911 580226 282920
rect 580172 282882 580224 282888
rect 580170 278896 580226 278905
rect 580170 278831 580226 278840
rect 580184 278798 580212 278831
rect 580172 278792 580224 278798
rect 580172 278734 580224 278740
rect 580170 274816 580226 274825
rect 580170 274751 580226 274760
rect 580184 274718 580212 274751
rect 580172 274712 580224 274718
rect 580172 274654 580224 274660
rect 579710 270736 579766 270745
rect 579710 270671 579766 270680
rect 579724 270570 579752 270671
rect 579712 270564 579764 270570
rect 579712 270506 579764 270512
rect 579618 266656 579674 266665
rect 579618 266591 579674 266600
rect 579632 266422 579660 266591
rect 579620 266416 579672 266422
rect 579620 266358 579672 266364
rect 580262 262576 580318 262585
rect 580262 262511 580318 262520
rect 580276 262274 580304 262511
rect 580264 262268 580316 262274
rect 580264 262210 580316 262216
rect 580262 258496 580318 258505
rect 580262 258431 580318 258440
rect 579802 254416 579858 254425
rect 579802 254351 579858 254360
rect 579816 253978 579844 254351
rect 579804 253972 579856 253978
rect 579804 253914 579856 253920
rect 579988 251184 580040 251190
rect 579988 251126 580040 251132
rect 580000 250345 580028 251126
rect 579986 250336 580042 250345
rect 579986 250271 580042 250280
rect 580170 242176 580226 242185
rect 580170 242111 580226 242120
rect 580184 241534 580212 242111
rect 580172 241528 580224 241534
rect 580172 241470 580224 241476
rect 580172 238740 580224 238746
rect 580172 238682 580224 238688
rect 580184 238105 580212 238682
rect 580170 238096 580226 238105
rect 580170 238031 580226 238040
rect 579986 225856 580042 225865
rect 579986 225791 580042 225800
rect 580000 225010 580028 225791
rect 579988 225004 580040 225010
rect 579988 224946 580040 224952
rect 580170 197976 580226 197985
rect 580170 197911 580226 197920
rect 580184 197402 580212 197911
rect 580172 197396 580224 197402
rect 580172 197338 580224 197344
rect 580276 197305 580304 258431
rect 580368 199345 580396 605231
rect 580538 588976 580594 588985
rect 580538 588911 580594 588920
rect 580446 379536 580502 379545
rect 580446 379471 580502 379480
rect 580354 199336 580410 199345
rect 580354 199271 580410 199280
rect 580262 197296 580318 197305
rect 580262 197231 580318 197240
rect 580356 196036 580408 196042
rect 580356 195978 580408 195984
rect 580264 194608 580316 194614
rect 580264 194550 580316 194556
rect 579802 193896 579858 193905
rect 579802 193831 579858 193840
rect 579816 193594 579844 193831
rect 579804 193588 579856 193594
rect 579804 193530 579856 193536
rect 579160 191820 579212 191826
rect 579160 191762 579212 191768
rect 579618 189816 579674 189825
rect 579068 189780 579120 189786
rect 579618 189751 579674 189760
rect 579068 189722 579120 189728
rect 579632 189106 579660 189751
rect 579620 189100 579672 189106
rect 579620 189042 579672 189048
rect 580276 185745 580304 194550
rect 580262 185736 580318 185745
rect 580262 185671 580318 185680
rect 580172 182096 580224 182102
rect 580172 182038 580224 182044
rect 580184 181665 580212 182038
rect 580170 181656 580226 181665
rect 580170 181591 580226 181600
rect 578976 179308 579028 179314
rect 578976 179250 579028 179256
rect 573362 178735 573418 178744
rect 577780 178764 577832 178770
rect 577780 178706 577832 178712
rect 560944 178696 560996 178702
rect 560944 178638 560996 178644
rect 580172 177880 580224 177886
rect 580172 177822 580224 177828
rect 580184 177585 580212 177822
rect 580170 177576 580226 177585
rect 580170 177511 580226 177520
rect 558274 176488 558330 176497
rect 558274 176423 558330 176432
rect 544382 176352 544438 176361
rect 544382 176287 544438 176296
rect 382278 176216 382334 176225
rect 382278 176151 382334 176160
rect 367098 176080 367154 176089
rect 367098 176015 367154 176024
rect 351918 175944 351974 175953
rect 351918 175879 351974 175888
rect 580170 173496 580226 173505
rect 580170 173431 580226 173440
rect 580184 173194 580212 173431
rect 580172 173188 580224 173194
rect 580172 173130 580224 173136
rect 580262 169416 580318 169425
rect 580262 169351 580318 169360
rect 580170 165336 580226 165345
rect 580170 165271 580226 165280
rect 580184 164286 580212 165271
rect 580172 164280 580224 164286
rect 580172 164222 580224 164228
rect 580170 161936 580226 161945
rect 580170 161871 580226 161880
rect 580184 161498 580212 161871
rect 580172 161492 580224 161498
rect 580172 161434 580224 161440
rect 579618 153776 579674 153785
rect 579618 153711 579674 153720
rect 579632 153270 579660 153711
rect 579620 153264 579672 153270
rect 579620 153206 579672 153212
rect 580172 149728 580224 149734
rect 580170 149696 580172 149705
rect 580224 149696 580226 149705
rect 580170 149631 580226 149640
rect 580172 146940 580224 146946
rect 580172 146882 580224 146888
rect 580184 145625 580212 146882
rect 580170 145616 580226 145625
rect 580170 145551 580226 145560
rect 580276 144906 580304 169351
rect 580264 144900 580316 144906
rect 580264 144842 580316 144848
rect 534080 143676 534132 143682
rect 534080 143618 534132 143624
rect 492680 143608 492732 143614
rect 492680 143550 492732 143556
rect 270500 142996 270552 143002
rect 270500 142938 270552 142944
rect 220820 142384 220872 142390
rect 220820 142326 220872 142332
rect 219808 66224 219860 66230
rect 219808 66166 219860 66172
rect 219716 60716 219768 60722
rect 219716 60658 219768 60664
rect 220728 60716 220780 60722
rect 220728 60658 220780 60664
rect 220740 60110 220768 60658
rect 220728 60104 220780 60110
rect 220728 60046 220780 60052
rect 219624 52420 219676 52426
rect 219624 52362 219676 52368
rect 220728 52420 220780 52426
rect 220728 52362 220780 52368
rect 220740 51746 220768 52362
rect 220728 51740 220780 51746
rect 220728 51682 220780 51688
rect 220832 16574 220860 142326
rect 255320 72480 255372 72486
rect 255320 72422 255372 72428
rect 236000 66972 236052 66978
rect 236000 66914 236052 66920
rect 231860 57316 231912 57322
rect 231860 57258 231912 57264
rect 224960 54596 225012 54602
rect 224960 54538 225012 54544
rect 216692 16546 217272 16574
rect 220832 16546 221136 16574
rect 211804 3052 211856 3058
rect 211804 2994 211856 3000
rect 213828 3052 213880 3058
rect 213828 2994 213880 3000
rect 213840 480 213868 2994
rect 206070 354 206182 480
rect 205652 326 206182 354
rect 202206 -960 202318 326
rect 206070 -960 206182 326
rect 209934 -960 210046 480
rect 213798 -960 213910 480
rect 217244 354 217272 16546
rect 217662 354 217774 480
rect 217244 326 217774 354
rect 221108 354 221136 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 224972 354 225000 54538
rect 231872 16574 231900 57258
rect 236012 16574 236040 66914
rect 251180 58744 251232 58750
rect 251180 58686 251232 58692
rect 242900 42152 242952 42158
rect 242900 42094 242952 42100
rect 231872 16546 232544 16574
rect 236012 16546 236408 16574
rect 232516 480 232544 16546
rect 236380 480 236408 16546
rect 242912 3602 242940 42094
rect 247040 35284 247092 35290
rect 247040 35226 247092 35232
rect 247052 16574 247080 35226
rect 251192 16574 251220 58686
rect 255332 16574 255360 72422
rect 265624 71120 265676 71126
rect 265624 71062 265676 71068
rect 262220 25628 262272 25634
rect 262220 25570 262272 25576
rect 247052 16546 248000 16574
rect 251192 16546 251864 16574
rect 255332 16546 255728 16574
rect 242900 3596 242952 3602
rect 242900 3538 242952 3544
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 244108 480 244136 3538
rect 247972 480 248000 16546
rect 251836 480 251864 16546
rect 255700 480 255728 16546
rect 262232 3602 262260 25570
rect 265636 3602 265664 71062
rect 270512 16574 270540 142938
rect 426440 142656 426492 142662
rect 426440 142598 426492 142604
rect 365720 142316 365772 142322
rect 365720 142258 365772 142264
rect 335360 140072 335412 140078
rect 335360 140014 335412 140020
rect 289820 76560 289872 76566
rect 289820 76502 289872 76508
rect 281540 75268 281592 75274
rect 281540 75210 281592 75216
rect 274640 73840 274692 73846
rect 274640 73782 274692 73788
rect 274652 16574 274680 73782
rect 278780 64252 278832 64258
rect 278780 64194 278832 64200
rect 278792 16574 278820 64194
rect 270512 16546 271184 16574
rect 274652 16546 275048 16574
rect 278792 16546 278912 16574
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 265624 3596 265676 3602
rect 265624 3538 265676 3544
rect 267280 3596 267332 3602
rect 267280 3538 267332 3544
rect 263428 480 263456 3538
rect 267292 480 267320 3538
rect 271156 480 271184 16546
rect 275020 480 275048 16546
rect 278884 480 278912 16546
rect 281552 3602 281580 75210
rect 281540 3596 281592 3602
rect 281540 3538 281592 3544
rect 282736 3596 282788 3602
rect 282736 3538 282788 3544
rect 282748 480 282776 3538
rect 289832 480 289860 76502
rect 300860 69760 300912 69766
rect 300860 69702 300912 69708
rect 296720 28348 296772 28354
rect 296720 28290 296772 28296
rect 296732 16574 296760 28290
rect 300872 16574 300900 69702
rect 309140 51808 309192 51814
rect 309140 51750 309192 51756
rect 305000 50448 305052 50454
rect 305000 50390 305052 50396
rect 296732 16546 297128 16574
rect 300872 16546 300992 16574
rect 225390 354 225502 480
rect 224972 326 225502 354
rect 217662 -960 217774 326
rect 221526 -960 221638 326
rect 225390 -960 225502 326
rect 228610 -960 228722 480
rect 232474 -960 232586 480
rect 236338 -960 236450 480
rect 240202 -960 240314 480
rect 244066 -960 244178 480
rect 247930 -960 248042 480
rect 251794 -960 251906 480
rect 255658 -960 255770 480
rect 259522 -960 259634 480
rect 263386 -960 263498 480
rect 267250 -960 267362 480
rect 271114 -960 271226 480
rect 274978 -960 275090 480
rect 278842 -960 278954 480
rect 282706 -960 282818 480
rect 285926 -960 286038 480
rect 289790 -960 289902 480
rect 293654 -960 293766 480
rect 297100 354 297128 16546
rect 297518 354 297630 480
rect 297100 326 297630 354
rect 300964 354 300992 16546
rect 301382 354 301494 480
rect 300964 326 301494 354
rect 305012 354 305040 50390
rect 309152 480 309180 51750
rect 324320 46232 324372 46238
rect 324320 46174 324372 46180
rect 320180 21480 320232 21486
rect 320180 21422 320232 21428
rect 320192 16574 320220 21422
rect 320192 16546 320312 16574
rect 316408 14544 316460 14550
rect 316408 14486 316460 14492
rect 305246 354 305358 480
rect 305012 326 305358 354
rect 297518 -960 297630 326
rect 301382 -960 301494 326
rect 305246 -960 305358 326
rect 309110 -960 309222 480
rect 312974 -960 313086 480
rect 316420 354 316448 14486
rect 316838 354 316950 480
rect 316420 326 316950 354
rect 320284 354 320312 16546
rect 320702 354 320814 480
rect 320284 326 320814 354
rect 324332 354 324360 46174
rect 331220 38004 331272 38010
rect 331220 37946 331272 37952
rect 331232 16574 331260 37946
rect 335372 16574 335400 140014
rect 346400 66292 346452 66298
rect 346400 66234 346452 66240
rect 342260 60036 342312 60042
rect 342260 59978 342312 59984
rect 342272 16574 342300 59978
rect 346412 16574 346440 66234
rect 354680 43512 354732 43518
rect 354680 43454 354732 43460
rect 350540 22840 350592 22846
rect 350540 22782 350592 22788
rect 350552 16574 350580 22782
rect 354692 16574 354720 43454
rect 357440 29708 357492 29714
rect 357440 29650 357492 29656
rect 331232 16546 331904 16574
rect 335372 16546 335768 16574
rect 342272 16546 343312 16574
rect 346412 16546 347176 16574
rect 350552 16546 351040 16574
rect 354692 16546 354904 16574
rect 324566 354 324678 480
rect 324332 326 324678 354
rect 316838 -960 316950 326
rect 320702 -960 320814 326
rect 324566 -960 324678 326
rect 328430 -960 328542 480
rect 331876 354 331904 16546
rect 332294 354 332406 480
rect 331876 326 332406 354
rect 335740 354 335768 16546
rect 340052 9036 340104 9042
rect 340052 8978 340104 8984
rect 340064 480 340092 8978
rect 343284 480 343312 16546
rect 347148 480 347176 16546
rect 351012 480 351040 16546
rect 354876 480 354904 16546
rect 357452 3602 357480 29650
rect 361580 18692 361632 18698
rect 361580 18634 361632 18640
rect 361592 16574 361620 18634
rect 365732 16574 365760 142258
rect 395344 141500 395396 141506
rect 395344 141442 395396 141448
rect 385040 61464 385092 61470
rect 385040 61406 385092 61412
rect 376760 55956 376812 55962
rect 376760 55898 376812 55904
rect 374000 49020 374052 49026
rect 374000 48962 374052 48968
rect 369860 47660 369912 47666
rect 369860 47602 369912 47608
rect 369872 16574 369900 47602
rect 374012 16574 374040 48962
rect 361592 16546 362632 16574
rect 365732 16546 366496 16574
rect 369872 16546 370360 16574
rect 374012 16546 374224 16574
rect 357440 3596 357492 3602
rect 357440 3538 357492 3544
rect 358728 3596 358780 3602
rect 358728 3538 358780 3544
rect 358740 480 358768 3538
rect 362604 480 362632 16546
rect 366468 480 366496 16546
rect 370332 480 370360 16546
rect 374196 480 374224 16546
rect 376772 2650 376800 55898
rect 385052 16574 385080 61406
rect 389180 37936 389232 37942
rect 389180 37878 389232 37884
rect 389192 16574 389220 37878
rect 392584 22772 392636 22778
rect 392584 22714 392636 22720
rect 385052 16546 385816 16574
rect 389192 16546 389680 16574
rect 381912 3528 381964 3534
rect 381912 3470 381964 3476
rect 376760 2644 376812 2650
rect 376760 2586 376812 2592
rect 378048 2644 378100 2650
rect 378048 2586 378100 2592
rect 378060 480 378088 2586
rect 381924 480 381952 3470
rect 385788 480 385816 16546
rect 389652 480 389680 16546
rect 392596 3058 392624 22714
rect 395356 3534 395384 141442
rect 407120 69692 407172 69698
rect 407120 69634 407172 69640
rect 404360 60104 404412 60110
rect 404360 60046 404412 60052
rect 400220 54528 400272 54534
rect 400220 54470 400272 54476
rect 396080 46300 396132 46306
rect 396080 46242 396132 46248
rect 395344 3528 395396 3534
rect 395344 3470 395396 3476
rect 392584 3052 392636 3058
rect 392584 2994 392636 3000
rect 393504 3052 393556 3058
rect 393504 2994 393556 3000
rect 393516 480 393544 2994
rect 396092 2650 396120 46242
rect 396080 2644 396132 2650
rect 396080 2586 396132 2592
rect 397368 2644 397420 2650
rect 397368 2586 397420 2592
rect 397380 480 397408 2586
rect 336158 354 336270 480
rect 335740 326 336270 354
rect 332294 -960 332406 326
rect 336158 -960 336270 326
rect 340022 -960 340134 480
rect 343242 -960 343354 480
rect 347106 -960 347218 480
rect 350970 -960 351082 480
rect 354834 -960 354946 480
rect 358698 -960 358810 480
rect 362562 -960 362674 480
rect 366426 -960 366538 480
rect 370290 -960 370402 480
rect 374154 -960 374266 480
rect 378018 -960 378130 480
rect 381882 -960 381994 480
rect 385746 -960 385858 480
rect 389610 -960 389722 480
rect 393474 -960 393586 480
rect 397338 -960 397450 480
rect 400232 354 400260 54470
rect 404372 16574 404400 60046
rect 407132 16574 407160 69634
rect 423680 33788 423732 33794
rect 423680 33730 423732 33736
rect 423692 16574 423720 33730
rect 426452 16574 426480 142598
rect 484400 71052 484452 71058
rect 484400 70994 484452 71000
rect 438860 65544 438912 65550
rect 438860 65486 438912 65492
rect 430580 62824 430632 62830
rect 430580 62766 430632 62772
rect 430592 16574 430620 62766
rect 434720 21412 434772 21418
rect 434720 21354 434772 21360
rect 434732 16574 434760 21354
rect 404372 16546 404492 16574
rect 407132 16546 407896 16574
rect 423692 16546 423812 16574
rect 426452 16546 427216 16574
rect 430592 16546 431080 16574
rect 434732 16546 434944 16574
rect 404464 480 404492 16546
rect 400558 354 400670 480
rect 400232 326 400670 354
rect 400558 -960 400670 326
rect 404422 -960 404534 480
rect 407868 354 407896 16546
rect 418804 10328 418856 10334
rect 418804 10270 418856 10276
rect 418816 3534 418844 10270
rect 416044 3528 416096 3534
rect 416044 3470 416096 3476
rect 418804 3528 418856 3534
rect 418804 3470 418856 3476
rect 419908 3528 419960 3534
rect 419908 3470 419960 3476
rect 416056 480 416084 3470
rect 419920 480 419948 3470
rect 423784 480 423812 16546
rect 408286 354 408398 480
rect 407868 326 408398 354
rect 408286 -960 408398 326
rect 412150 -960 412262 480
rect 416014 -960 416126 480
rect 419878 -960 419990 480
rect 423742 -960 423854 480
rect 427188 354 427216 16546
rect 427606 354 427718 480
rect 427188 326 427718 354
rect 431052 354 431080 16546
rect 431470 354 431582 480
rect 431052 326 431582 354
rect 434916 354 434944 16546
rect 435334 354 435446 480
rect 434916 326 435446 354
rect 438872 354 438900 65486
rect 469220 53100 469272 53106
rect 469220 53042 469272 53048
rect 442264 47592 442316 47598
rect 442264 47534 442316 47540
rect 442276 3534 442304 47534
rect 456800 43444 456852 43450
rect 456800 43386 456852 43392
rect 454040 18624 454092 18630
rect 454040 18566 454092 18572
rect 454052 16574 454080 18566
rect 456812 16574 456840 43386
rect 465080 17264 465132 17270
rect 465080 17206 465132 17212
rect 465092 16574 465120 17206
rect 469232 16574 469260 53042
rect 480260 26920 480312 26926
rect 480260 26862 480312 26868
rect 480272 16574 480300 26862
rect 484412 16574 484440 70994
rect 488540 64184 488592 64190
rect 488540 64126 488592 64132
rect 488552 16574 488580 64126
rect 454052 16546 454264 16574
rect 456812 16546 457944 16574
rect 465092 16546 465672 16574
rect 469232 16546 469536 16574
rect 480272 16546 481128 16574
rect 484412 16546 484992 16574
rect 488552 16546 488856 16574
rect 442264 3528 442316 3534
rect 442264 3470 442316 3476
rect 443092 3528 443144 3534
rect 443092 3470 443144 3476
rect 443104 480 443132 3470
rect 439198 354 439310 480
rect 438872 326 439310 354
rect 427606 -960 427718 326
rect 431470 -960 431582 326
rect 435334 -960 435446 326
rect 439198 -960 439310 326
rect 443062 -960 443174 480
rect 446926 -960 447038 480
rect 450790 -960 450902 480
rect 454236 354 454264 16546
rect 457916 480 457944 16546
rect 461768 7608 461820 7614
rect 461768 7550 461820 7556
rect 461780 480 461808 7550
rect 465644 480 465672 16546
rect 469508 480 469536 16546
rect 477224 13116 477276 13122
rect 477224 13058 477276 13064
rect 473360 6180 473412 6186
rect 473360 6122 473412 6128
rect 473372 480 473400 6122
rect 477236 480 477264 13058
rect 481100 480 481128 16546
rect 484964 480 484992 16546
rect 488828 480 488856 16546
rect 492692 480 492720 143550
rect 514760 142588 514812 142594
rect 514760 142530 514812 142536
rect 503720 66904 503772 66910
rect 503720 66846 503772 66852
rect 499580 35216 499632 35222
rect 499580 35158 499632 35164
rect 495440 31068 495492 31074
rect 495440 31010 495492 31016
rect 495452 16574 495480 31010
rect 499592 16574 499620 35158
rect 503732 16574 503760 66846
rect 510620 58676 510672 58682
rect 510620 58618 510672 58624
rect 507860 29640 507912 29646
rect 507860 29582 507912 29588
rect 507872 16574 507900 29582
rect 510632 16574 510660 58618
rect 495452 16546 496584 16574
rect 499592 16546 500448 16574
rect 503732 16546 504312 16574
rect 507872 16546 508176 16574
rect 510632 16546 510936 16574
rect 496556 480 496584 16546
rect 500420 480 500448 16546
rect 504284 480 504312 16546
rect 508148 480 508176 16546
rect 454654 354 454766 480
rect 454236 326 454766 354
rect 454654 -960 454766 326
rect 457874 -960 457986 480
rect 461738 -960 461850 480
rect 465602 -960 465714 480
rect 469466 -960 469578 480
rect 473330 -960 473442 480
rect 477194 -960 477306 480
rect 481058 -960 481170 480
rect 484922 -960 485034 480
rect 488786 -960 488898 480
rect 492650 -960 492762 480
rect 496514 -960 496626 480
rect 500378 -960 500490 480
rect 504242 -960 504354 480
rect 508106 -960 508218 480
rect 510908 354 510936 16546
rect 511326 354 511438 480
rect 510908 326 511438 354
rect 514772 354 514800 142530
rect 518900 141432 518952 141438
rect 518900 141374 518952 141380
rect 515190 354 515302 480
rect 514772 326 515302 354
rect 518912 354 518940 141374
rect 525800 75200 525852 75206
rect 525800 75142 525852 75148
rect 521660 42084 521712 42090
rect 521660 42026 521712 42032
rect 521672 16574 521700 42026
rect 525812 16574 525840 75142
rect 521672 16546 522528 16574
rect 525812 16546 526392 16574
rect 519054 354 519166 480
rect 518912 326 519166 354
rect 522500 354 522528 16546
rect 522918 354 523030 480
rect 522500 326 523030 354
rect 526364 354 526392 16546
rect 530676 8968 530728 8974
rect 530676 8910 530728 8916
rect 530688 480 530716 8910
rect 526782 354 526894 480
rect 526364 326 526894 354
rect 511326 -960 511438 326
rect 515190 -960 515302 326
rect 519054 -960 519166 326
rect 522918 -960 523030 326
rect 526782 -960 526894 326
rect 530646 -960 530758 480
rect 534092 354 534120 143618
rect 580264 142928 580316 142934
rect 580264 142870 580316 142876
rect 579618 142760 579674 142769
rect 579618 142695 579674 142704
rect 558184 61396 558236 61402
rect 558184 61338 558236 61344
rect 538220 55888 538272 55894
rect 538220 55830 538272 55836
rect 534510 354 534622 480
rect 534092 326 534622 354
rect 538232 354 538260 55830
rect 543004 50380 543056 50386
rect 543004 50322 543056 50328
rect 543016 5506 543044 50322
rect 549536 14476 549588 14482
rect 549536 14418 549588 14424
rect 543004 5500 543056 5506
rect 543004 5442 543056 5448
rect 542268 4820 542320 4826
rect 542268 4762 542320 4768
rect 542280 480 542308 4762
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 534510 -960 534622 326
rect 538374 -960 538486 326
rect 542238 -960 542350 480
rect 546102 -960 546214 480
rect 549548 354 549576 14418
rect 558196 3466 558224 61338
rect 560300 57248 560352 57254
rect 560300 57190 560352 57196
rect 560312 16574 560340 57190
rect 563704 51740 563756 51746
rect 563704 51682 563756 51688
rect 560312 16546 561168 16574
rect 557724 3460 557776 3466
rect 557724 3402 557776 3408
rect 558184 3460 558236 3466
rect 558184 3402 558236 3408
rect 557736 480 557764 3402
rect 549966 354 550078 480
rect 549548 326 550078 354
rect 549966 -960 550078 326
rect 553830 -960 553942 480
rect 557694 -960 557806 480
rect 561140 354 561168 16546
rect 563716 3058 563744 51682
rect 578884 39364 578936 39370
rect 578884 39306 578936 39312
rect 571340 28280 571392 28286
rect 571340 28222 571392 28228
rect 571352 3534 571380 28222
rect 575480 25560 575532 25566
rect 575480 25502 575532 25508
rect 575492 16574 575520 25502
rect 575492 16546 576440 16574
rect 571340 3528 571392 3534
rect 571340 3470 571392 3476
rect 572536 3528 572588 3534
rect 572536 3470 572588 3476
rect 568672 3460 568724 3466
rect 568672 3402 568724 3408
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 565452 3052 565504 3058
rect 565452 2994 565504 3000
rect 565464 480 565492 2994
rect 568684 480 568712 3402
rect 572548 480 572576 3470
rect 576412 480 576440 16546
rect 561558 354 561670 480
rect 561140 326 561670 354
rect 561558 -960 561670 326
rect 565422 -960 565534 480
rect 568642 -960 568754 480
rect 572506 -960 572618 480
rect 576370 -960 576482 480
rect 578896 105 578924 39306
rect 579632 6914 579660 142695
rect 580170 137456 580226 137465
rect 580170 137391 580226 137400
rect 580184 136678 580212 137391
rect 580172 136672 580224 136678
rect 580172 136614 580224 136620
rect 580170 125216 580226 125225
rect 580170 125151 580226 125160
rect 580184 124234 580212 125151
rect 580172 124228 580224 124234
rect 580172 124170 580224 124176
rect 580170 112976 580226 112985
rect 580170 112911 580226 112920
rect 580184 112470 580212 112911
rect 580172 112464 580224 112470
rect 580172 112406 580224 112412
rect 580170 85096 580226 85105
rect 580170 85031 580226 85040
rect 580184 80034 580212 85031
rect 580172 80028 580224 80034
rect 580172 79970 580224 79976
rect 580276 72865 580304 142870
rect 580368 129305 580396 195978
rect 580460 193186 580488 379471
rect 580552 199481 580580 588911
rect 580630 327176 580686 327185
rect 580630 327111 580686 327120
rect 580538 199472 580594 199481
rect 580538 199407 580594 199416
rect 580644 193934 580672 327111
rect 580722 229936 580778 229945
rect 580722 229871 580778 229880
rect 580736 200802 580764 229871
rect 580814 214296 580870 214305
rect 580814 214231 580870 214240
rect 580724 200796 580776 200802
rect 580724 200738 580776 200744
rect 580828 195294 580856 214231
rect 580906 210216 580962 210225
rect 580906 210151 580962 210160
rect 580816 195288 580868 195294
rect 580816 195230 580868 195236
rect 580632 193928 580684 193934
rect 580632 193870 580684 193876
rect 580448 193180 580500 193186
rect 580448 193122 580500 193128
rect 580920 192574 580948 210151
rect 580908 192568 580960 192574
rect 580908 192510 580960 192516
rect 581012 185609 581040 703582
rect 582024 703474 582052 703582
rect 582166 703520 582278 704960
rect 582208 703474 582236 703520
rect 582024 703446 582236 703474
rect 582378 690296 582434 690305
rect 582378 690231 582434 690240
rect 581734 661736 581790 661745
rect 581734 661671 581790 661680
rect 581642 657656 581698 657665
rect 581642 657591 581698 657600
rect 580998 185600 581054 185609
rect 580998 185535 581054 185544
rect 581656 179382 581684 657591
rect 581748 194041 581776 661671
rect 581826 440056 581882 440065
rect 581826 439991 581882 440000
rect 581734 194032 581790 194041
rect 581734 193967 581790 193976
rect 581840 184890 581868 439991
rect 581828 184884 581880 184890
rect 581828 184826 581880 184832
rect 582392 182918 582420 690231
rect 582470 682136 582526 682145
rect 582470 682071 582526 682080
rect 582380 182912 582432 182918
rect 582484 182889 582512 682071
rect 582654 637936 582710 637945
rect 582654 637871 582710 637880
rect 582562 621616 582618 621625
rect 582562 621551 582618 621560
rect 582576 183161 582604 621551
rect 582668 200705 582696 637871
rect 582838 617536 582894 617545
rect 582838 617471 582894 617480
rect 582746 613456 582802 613465
rect 582746 613391 582802 613400
rect 582654 200696 582710 200705
rect 582654 200631 582710 200640
rect 582760 190466 582788 613391
rect 582852 195537 582880 617471
rect 582930 557016 582986 557025
rect 582930 556951 582986 556960
rect 582838 195528 582894 195537
rect 582838 195463 582894 195472
rect 582748 190460 582800 190466
rect 582748 190402 582800 190408
rect 582562 183152 582618 183161
rect 582562 183087 582618 183096
rect 582380 182854 582432 182860
rect 582470 182880 582526 182889
rect 582470 182815 582526 182824
rect 582944 180713 582972 556951
rect 583022 532536 583078 532545
rect 583022 532471 583078 532480
rect 583036 182850 583064 532471
rect 583024 182844 583076 182850
rect 583024 182786 583076 182792
rect 582930 180704 582986 180713
rect 582930 180639 582986 180648
rect 581644 179376 581696 179382
rect 581644 179318 581696 179324
rect 580538 147792 580594 147801
rect 580538 147727 580594 147736
rect 580448 146328 580500 146334
rect 580448 146270 580500 146276
rect 580460 141545 580488 146270
rect 580446 141536 580502 141545
rect 580446 141471 580502 141480
rect 580448 139460 580500 139466
rect 580448 139402 580500 139408
rect 580354 129296 580410 129305
rect 580354 129231 580410 129240
rect 580460 108905 580488 139402
rect 580552 117065 580580 147727
rect 580724 142860 580776 142866
rect 580724 142802 580776 142808
rect 580632 138712 580684 138718
rect 580632 138654 580684 138660
rect 580644 121145 580672 138654
rect 580736 133385 580764 142802
rect 580722 133376 580778 133385
rect 580722 133311 580778 133320
rect 580630 121136 580686 121145
rect 580630 121071 580686 121080
rect 580538 117056 580594 117065
rect 580538 116991 580594 117000
rect 580446 108896 580502 108905
rect 580446 108831 580502 108840
rect 580354 104816 580410 104825
rect 580354 104751 580410 104760
rect 580262 72856 580318 72865
rect 580262 72791 580318 72800
rect 579988 69012 580040 69018
rect 579988 68954 580040 68960
rect 580000 68785 580028 68954
rect 579986 68776 580042 68785
rect 579986 68711 580042 68720
rect 580368 63510 580396 104751
rect 580630 101416 580686 101425
rect 580630 101351 580686 101360
rect 580446 97336 580502 97345
rect 580446 97271 580502 97280
rect 580356 63504 580408 63510
rect 580356 63446 580408 63452
rect 580460 62121 580488 97271
rect 580538 89176 580594 89185
rect 580538 89111 580594 89120
rect 580552 63442 580580 89111
rect 580644 79762 580672 101351
rect 580722 93256 580778 93265
rect 580722 93191 580778 93200
rect 580632 79756 580684 79762
rect 580632 79698 580684 79704
rect 580630 76936 580686 76945
rect 580630 76871 580686 76880
rect 580644 67590 580672 76871
rect 580736 72321 580764 93191
rect 580722 72312 580778 72321
rect 580722 72247 580778 72256
rect 580632 67584 580684 67590
rect 580632 67526 580684 67532
rect 580540 63436 580592 63442
rect 580540 63378 580592 63384
rect 580446 62112 580502 62121
rect 580446 62047 580502 62056
rect 580172 49700 580224 49706
rect 580172 49642 580224 49648
rect 580184 48385 580212 49642
rect 580170 48376 580226 48385
rect 580170 48311 580226 48320
rect 579988 45552 580040 45558
rect 579988 45494 580040 45500
rect 580000 44305 580028 45494
rect 579986 44296 580042 44305
rect 579986 44231 580042 44240
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 40905 580212 41346
rect 580170 40896 580226 40905
rect 580170 40831 580226 40840
rect 580172 37256 580224 37262
rect 580172 37198 580224 37204
rect 580184 36825 580212 37198
rect 580170 36816 580226 36825
rect 580170 36751 580226 36760
rect 580172 33108 580224 33114
rect 580172 33050 580224 33056
rect 580184 32745 580212 33050
rect 580170 32736 580226 32745
rect 580170 32671 580226 32680
rect 580172 24812 580224 24818
rect 580172 24754 580224 24760
rect 580184 24585 580212 24754
rect 580170 24576 580226 24585
rect 580170 24511 580226 24520
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 20505 580212 20606
rect 580170 20496 580226 20505
rect 580170 20431 580226 20440
rect 580172 16584 580224 16590
rect 580172 16526 580224 16532
rect 580184 16425 580212 16526
rect 580170 16416 580226 16425
rect 580170 16351 580226 16360
rect 580172 12436 580224 12442
rect 580172 12378 580224 12384
rect 580184 12345 580212 12378
rect 580170 12336 580226 12345
rect 580170 12271 580226 12280
rect 580172 8288 580224 8294
rect 580170 8256 580172 8265
rect 580224 8256 580226 8265
rect 580170 8191 580226 8200
rect 579632 6886 580304 6914
rect 580172 5500 580224 5506
rect 580172 5442 580224 5448
rect 580184 4185 580212 5442
rect 580170 4176 580226 4185
rect 580170 4111 580226 4120
rect 580276 480 580304 6886
rect 578882 96 578938 105
rect 578882 31 578938 40
rect 580234 -960 580346 480
<< via2 >>
rect 3054 701800 3110 701856
rect 3146 693640 3202 693696
rect 3422 689560 3478 689616
rect 3146 685480 3202 685536
rect 3422 681400 3478 681456
rect 3238 673240 3294 673296
rect 3422 669160 3478 669216
rect 3238 665080 3294 665136
rect 3422 661036 3424 661056
rect 3424 661036 3476 661056
rect 3476 661036 3478 661056
rect 3422 661000 3478 661036
rect 3054 653520 3110 653576
rect 3422 645360 3478 645416
rect 3422 629040 3478 629096
rect 3238 624960 3294 625016
rect 3422 620880 3478 620936
rect 3238 616800 3294 616856
rect 3422 612756 3424 612776
rect 3424 612756 3476 612776
rect 3476 612756 3478 612776
rect 3422 612720 3478 612756
rect 3422 608660 3478 608696
rect 3422 608640 3424 608660
rect 3424 608640 3476 608660
rect 3476 608640 3478 608660
rect 3422 604560 3478 604616
rect 3422 600480 3478 600536
rect 3422 597080 3478 597136
rect 3422 588920 3478 588976
rect 3422 584840 3478 584896
rect 3422 580760 3478 580816
rect 3238 576680 3294 576736
rect 3422 572600 3478 572656
rect 3238 568520 3294 568576
rect 3422 564460 3478 564496
rect 3422 564440 3424 564460
rect 3424 564440 3476 564460
rect 3476 564440 3478 564460
rect 3422 560360 3478 560416
rect 3422 556280 3478 556336
rect 3422 552200 3478 552256
rect 3238 548120 3294 548176
rect 3330 544040 3386 544096
rect 3422 539960 3478 540016
rect 3238 532480 3294 532536
rect 3422 528400 3478 528456
rect 3238 524320 3294 524376
rect 3422 520276 3424 520296
rect 3424 520276 3476 520296
rect 3476 520276 3478 520296
rect 3422 520240 3478 520276
rect 3422 516180 3478 516216
rect 3422 516160 3424 516180
rect 3424 516160 3476 516180
rect 3476 516160 3478 516180
rect 3422 512080 3478 512136
rect 3422 508000 3478 508056
rect 3238 503920 3294 503976
rect 3330 499840 3386 499896
rect 2870 495760 2926 495816
rect 3422 491680 3478 491736
rect 3422 487600 3478 487656
rect 3514 483520 3570 483576
rect 3422 480120 3478 480176
rect 3238 476040 3294 476096
rect 3422 471996 3424 472016
rect 3424 471996 3476 472016
rect 3476 471996 3478 472016
rect 3422 471960 3478 471996
rect 3422 467900 3478 467936
rect 3422 467880 3424 467900
rect 3424 467880 3476 467900
rect 3476 467880 3478 467900
rect 3422 463800 3478 463856
rect 3422 459720 3478 459776
rect 3238 455640 3294 455696
rect 3330 451560 3386 451616
rect 3422 443400 3478 443456
rect 3422 439320 3478 439376
rect 2870 427080 2926 427136
rect 2962 423000 3018 423056
rect 3330 403280 3386 403336
rect 2870 378800 2926 378856
rect 2962 374720 3018 374776
rect 3054 370640 3110 370696
rect 3054 362480 3110 362536
rect 3330 359080 3386 359136
rect 3330 355000 3386 355056
rect 3330 346840 3386 346896
rect 2962 330520 3018 330576
rect 3054 322360 3110 322416
rect 3054 314200 3110 314256
rect 3146 310120 3202 310176
rect 3238 306040 3294 306096
rect 3146 301960 3202 302016
rect 3330 298560 3386 298616
rect 2870 286320 2926 286376
rect 2962 282240 3018 282296
rect 3054 278160 3110 278216
rect 3054 270000 3110 270056
rect 3146 265920 3202 265976
rect 3054 261840 3110 261896
rect 3238 257760 3294 257816
rect 3146 253680 3202 253736
rect 3330 241440 3386 241496
rect 3330 229880 3386 229936
rect 3054 221720 3110 221776
rect 3146 209480 3202 209536
rect 3146 197240 3202 197296
rect 3514 431160 3570 431216
rect 3514 419600 3570 419656
rect 3514 415520 3570 415576
rect 3514 411440 3570 411496
rect 3514 407360 3570 407416
rect 3514 391040 3570 391096
rect 3514 386960 3570 387016
rect 3514 350920 3570 350976
rect 3514 342760 3570 342816
rect 3514 338680 3570 338736
rect 3514 318280 3570 318336
rect 3514 294480 3570 294536
rect 3514 290400 3570 290456
rect 3514 274080 3570 274136
rect 3514 249600 3570 249656
rect 3606 225800 3662 225856
rect 4066 201320 4122 201376
rect 4158 199280 4214 199336
rect 3422 193160 3478 193216
rect 3422 189100 3478 189136
rect 3422 189080 3424 189100
rect 3424 189080 3476 189100
rect 3476 189080 3478 189100
rect 3422 185000 3478 185056
rect 3422 180920 3478 180976
rect 3330 177520 3386 177576
rect 3422 173440 3478 173496
rect 3146 169360 3202 169416
rect 2778 165316 2780 165336
rect 2780 165316 2832 165336
rect 2832 165316 2834 165336
rect 2778 165280 2834 165316
rect 3514 161200 3570 161256
rect 3514 157120 3570 157176
rect 3514 153040 3570 153096
rect 3422 148996 3424 149016
rect 3424 148996 3476 149016
rect 3476 148996 3478 149016
rect 3422 148960 3478 148996
rect 3422 144916 3424 144936
rect 3424 144916 3476 144936
rect 3476 144916 3478 144936
rect 3422 144880 3478 144916
rect 31022 199416 31078 199472
rect 27618 193840 27674 193896
rect 38658 265512 38714 265568
rect 34518 193160 34574 193216
rect 12438 190168 12494 190224
rect 42798 187584 42854 187640
rect 62118 196968 62174 197024
rect 78034 200640 78090 200696
rect 77942 188264 77998 188320
rect 49698 186088 49754 186144
rect 88982 193976 89038 194032
rect 89074 190984 89130 191040
rect 92478 202136 92534 202192
rect 94502 188808 94558 188864
rect 3514 140800 3570 140856
rect 3422 136720 3478 136776
rect 3146 120400 3202 120456
rect 3238 117000 3294 117056
rect 3422 112920 3478 112976
rect 3422 108840 3478 108896
rect 3422 104760 3478 104816
rect 3330 100680 3386 100736
rect 3422 96636 3424 96656
rect 3424 96636 3476 96656
rect 3476 96636 3478 96656
rect 3422 96600 3478 96636
rect 3146 92520 3202 92576
rect 3422 84360 3478 84416
rect 3422 80280 3478 80336
rect 2778 76200 2834 76256
rect 3146 72120 3202 72176
rect 3146 68040 3202 68096
rect 3146 63960 3202 64016
rect 3422 56516 3424 56536
rect 3424 56516 3476 56536
rect 3476 56516 3478 56536
rect 3422 56480 3478 56516
rect 3422 52420 3478 52456
rect 3422 52400 3424 52420
rect 3424 52400 3476 52420
rect 3476 52400 3478 52420
rect 3238 48320 3294 48376
rect 3146 36080 3202 36136
rect 3146 32000 3202 32056
rect 3146 27920 3202 27976
rect 3054 23840 3110 23896
rect 3054 11600 3110 11656
rect 2962 7520 3018 7576
rect 3514 44240 3570 44296
rect 3514 40160 3570 40216
rect 3514 19760 3570 19816
rect 3514 15680 3570 15736
rect 3146 3440 3202 3496
rect 95054 200640 95110 200696
rect 95054 200096 95110 200152
rect 96342 195200 96398 195256
rect 97078 141752 97134 141808
rect 97078 75656 97134 75712
rect 96986 74976 97042 75032
rect 97630 191120 97686 191176
rect 98642 193024 98698 193080
rect 98826 188536 98882 188592
rect 97722 67496 97778 67552
rect 97630 64776 97686 64832
rect 98550 71032 98606 71088
rect 99010 81096 99066 81152
rect 99194 188264 99250 188320
rect 99194 74160 99250 74216
rect 98918 67224 98974 67280
rect 100206 81912 100262 81968
rect 100114 69808 100170 69864
rect 101494 80960 101550 81016
rect 101586 79056 101642 79112
rect 101678 77152 101734 77208
rect 102966 195744 103022 195800
rect 102690 81776 102746 81832
rect 102966 79464 103022 79520
rect 102874 78920 102930 78976
rect 104162 72664 104218 72720
rect 103334 64504 103390 64560
rect 104714 195336 104770 195392
rect 105634 200232 105690 200288
rect 105542 196832 105598 196888
rect 105818 79192 105874 79248
rect 105726 70896 105782 70952
rect 106922 191664 106978 191720
rect 107382 202136 107438 202192
rect 107382 201456 107438 201512
rect 107106 68312 107162 68368
rect 108210 139032 108266 139088
rect 108394 81232 108450 81288
rect 108210 76880 108266 76936
rect 108670 73888 108726 73944
rect 109038 188536 109094 188592
rect 109038 188264 109094 188320
rect 109498 78784 109554 78840
rect 109406 75384 109462 75440
rect 110142 188264 110198 188320
rect 110878 72800 110934 72856
rect 111154 83408 111210 83464
rect 111798 200640 111854 200696
rect 111890 191120 111946 191176
rect 114006 143112 114062 143168
rect 115202 138896 115258 138952
rect 115386 142704 115442 142760
rect 115386 140256 115442 140312
rect 114926 75520 114982 75576
rect 115846 138080 115902 138136
rect 115846 92520 115902 92576
rect 115846 81504 115902 81560
rect 116398 76200 116454 76256
rect 116582 145560 116638 145616
rect 117042 198872 117098 198928
rect 117134 139440 117190 139496
rect 116858 71168 116914 71224
rect 118146 71576 118202 71632
rect 118698 200912 118754 200968
rect 118698 199552 118754 199608
rect 118422 137944 118478 138000
rect 118514 73072 118570 73128
rect 119710 191120 119766 191176
rect 120630 218048 120686 218104
rect 119894 138624 119950 138680
rect 119802 75792 119858 75848
rect 119986 78512 120042 78568
rect 122562 262656 122618 262712
rect 121550 262248 121606 262304
rect 122562 259936 122618 259992
rect 129370 259664 129426 259720
rect 135442 263744 135498 263800
rect 136546 263744 136602 263800
rect 134890 262792 134946 262848
rect 138110 260072 138166 260128
rect 148046 263880 148102 263936
rect 131854 259528 131910 259584
rect 168930 263608 168986 263664
rect 179418 262792 179474 262848
rect 181442 262384 181498 262440
rect 183006 262928 183062 262984
rect 182178 259936 182234 259992
rect 183374 259936 183430 259992
rect 185490 262520 185546 262576
rect 184938 259936 184994 259992
rect 185858 259936 185914 259992
rect 183374 259528 183430 259584
rect 186962 259256 187018 259312
rect 122838 200640 122894 200696
rect 120722 180920 120778 180976
rect 120630 139032 120686 139088
rect 120722 138488 120778 138544
rect 121366 194520 121422 194576
rect 121734 122712 121790 122768
rect 121734 113192 121790 113248
rect 121734 113056 121790 113112
rect 121734 103536 121790 103592
rect 121734 103400 121790 103456
rect 121734 93880 121790 93936
rect 121734 93744 121790 93800
rect 123206 200368 123262 200424
rect 122838 197376 122894 197432
rect 122838 195880 122894 195936
rect 124126 198192 124182 198248
rect 124126 197376 124182 197432
rect 123482 193840 123538 193896
rect 124034 192480 124090 192536
rect 123482 179424 123538 179480
rect 124034 179424 124090 179480
rect 129002 200640 129058 200696
rect 127162 199824 127218 199880
rect 126150 199688 126206 199744
rect 125598 199008 125654 199064
rect 126886 198056 126942 198112
rect 124770 197648 124826 197704
rect 125506 197512 125562 197568
rect 125414 197104 125470 197160
rect 124770 179560 124826 179616
rect 124402 143112 124458 143168
rect 124310 139848 124366 139904
rect 127714 198464 127770 198520
rect 126978 194248 127034 194304
rect 125874 139576 125930 139632
rect 124126 139440 124182 139496
rect 127898 192480 127954 192536
rect 127714 179696 127770 179752
rect 126978 148552 127034 148608
rect 131486 200368 131542 200424
rect 131486 200096 131542 200152
rect 131670 200096 131726 200152
rect 131026 199824 131082 199880
rect 129002 197376 129058 197432
rect 128910 193840 128966 193896
rect 124034 139304 124090 139360
rect 125966 139304 126022 139360
rect 128450 139304 128506 139360
rect 132038 200252 132094 200288
rect 132038 200232 132040 200252
rect 132040 200232 132092 200252
rect 132092 200232 132094 200252
rect 132222 200232 132278 200288
rect 131854 199980 131910 200016
rect 131854 199960 131856 199980
rect 131856 199960 131908 199980
rect 131908 199960 131910 199980
rect 131854 199844 131910 199880
rect 131854 199824 131856 199844
rect 131856 199824 131908 199844
rect 131908 199824 131910 199844
rect 177946 200232 178002 200288
rect 132038 199824 132094 199880
rect 131946 199552 132002 199608
rect 131762 197940 131818 197976
rect 131762 197920 131764 197940
rect 131764 197920 131816 197940
rect 131816 197920 131818 197940
rect 131762 197240 131818 197296
rect 130566 195472 130622 195528
rect 130106 145968 130162 146024
rect 131854 197104 131910 197160
rect 130842 141888 130898 141944
rect 130474 140392 130530 140448
rect 132314 197240 132370 197296
rect 133188 199858 133244 199914
rect 132590 196424 132646 196480
rect 132406 196288 132462 196344
rect 133372 199824 133428 199880
rect 133142 199552 133198 199608
rect 132590 145832 132646 145888
rect 132130 140528 132186 140584
rect 133556 199858 133612 199914
rect 133832 199858 133888 199914
rect 134200 199824 134256 199880
rect 133602 199144 133658 199200
rect 133510 198328 133566 198384
rect 133510 197648 133566 197704
rect 133234 190440 133290 190496
rect 134384 199824 134440 199880
rect 134062 199552 134118 199608
rect 134752 199824 134808 199880
rect 134614 198192 134670 198248
rect 134338 193296 134394 193352
rect 134706 194248 134762 194304
rect 135120 199858 135176 199914
rect 134890 195608 134946 195664
rect 135074 196696 135130 196752
rect 135488 199824 135544 199880
rect 135672 199824 135728 199880
rect 135442 199688 135498 199744
rect 135258 197920 135314 197976
rect 135534 199552 135590 199608
rect 135948 199688 136004 199744
rect 136500 199824 136556 199880
rect 135902 198736 135958 198792
rect 136270 199144 136326 199200
rect 136178 195880 136234 195936
rect 136454 195880 136510 195936
rect 136868 199824 136924 199880
rect 136638 198192 136694 198248
rect 136638 197784 136694 197840
rect 136638 196016 136694 196072
rect 136822 199552 136878 199608
rect 136822 197784 136878 197840
rect 136822 197376 136878 197432
rect 136730 195880 136786 195936
rect 136638 195336 136694 195392
rect 137880 199824 137936 199880
rect 137098 198600 137154 198656
rect 137190 198464 137246 198520
rect 137374 196152 137430 196208
rect 136546 179424 136602 179480
rect 136454 177792 136510 177848
rect 136822 176160 136878 176216
rect 134522 141752 134578 141808
rect 136730 145696 136786 145752
rect 135994 142976 136050 143032
rect 137282 190304 137338 190360
rect 137282 179424 137338 179480
rect 138156 199824 138212 199880
rect 138432 199824 138488 199880
rect 137926 199552 137982 199608
rect 137834 199144 137890 199200
rect 138018 198464 138074 198520
rect 138294 198192 138350 198248
rect 138294 197512 138350 197568
rect 138202 196696 138258 196752
rect 138386 196152 138442 196208
rect 139076 199824 139132 199880
rect 139352 199824 139408 199880
rect 139536 199824 139592 199880
rect 138754 198192 138810 198248
rect 138386 195880 138442 195936
rect 137282 140664 137338 140720
rect 139030 199008 139086 199064
rect 138938 197376 138994 197432
rect 139122 195880 139178 195936
rect 139030 183504 139086 183560
rect 140088 199824 140144 199880
rect 140272 199824 140328 199880
rect 139306 199144 139362 199200
rect 139674 198056 139730 198112
rect 140226 199688 140282 199744
rect 140042 199552 140098 199608
rect 140042 199144 140098 199200
rect 141468 199824 141524 199880
rect 140502 196696 140558 196752
rect 141652 199824 141708 199880
rect 140962 198192 141018 198248
rect 140870 197784 140926 197840
rect 141238 196424 141294 196480
rect 141422 198736 141478 198792
rect 142112 199824 142168 199880
rect 142480 199824 142536 199880
rect 142940 199824 142996 199880
rect 142434 199724 142436 199744
rect 142436 199724 142488 199744
rect 142488 199724 142490 199744
rect 142434 199688 142490 199724
rect 143216 199824 143272 199880
rect 142342 199552 142398 199608
rect 142250 198464 142306 198520
rect 142158 198328 142214 198384
rect 141974 197104 142030 197160
rect 141422 177928 141478 177984
rect 140962 176432 141018 176488
rect 140870 176024 140926 176080
rect 142710 198736 142766 198792
rect 143078 199008 143134 199064
rect 142986 198736 143042 198792
rect 142526 180512 142582 180568
rect 142526 179968 142582 180024
rect 143262 199688 143318 199744
rect 143446 199552 143502 199608
rect 143354 196696 143410 196752
rect 143170 195880 143226 195936
rect 142986 195064 143042 195120
rect 144504 199824 144560 199880
rect 143446 188672 143502 188728
rect 142986 187040 143042 187096
rect 144090 199144 144146 199200
rect 143998 195472 144054 195528
rect 143446 182164 143502 182200
rect 143446 182144 143448 182164
rect 143448 182144 143500 182164
rect 143500 182144 143502 182164
rect 142802 148416 142858 148472
rect 144734 199552 144790 199608
rect 144366 197104 144422 197160
rect 144182 194520 144238 194576
rect 144182 183368 144238 183424
rect 144182 182688 144238 182744
rect 141514 140120 141570 140176
rect 144734 199008 144790 199064
rect 145792 199824 145848 199880
rect 145010 194520 145066 194576
rect 144642 188980 144644 189000
rect 144644 188980 144696 189000
rect 144696 188980 144698 189000
rect 144642 188944 144698 188980
rect 144734 186224 144790 186280
rect 144182 144336 144238 144392
rect 146436 199858 146492 199914
rect 146712 199858 146768 199914
rect 147080 199858 147136 199914
rect 147356 199858 147412 199914
rect 146850 199688 146906 199744
rect 146206 197648 146262 197704
rect 146114 197104 146170 197160
rect 146114 196560 146170 196616
rect 146574 199572 146630 199608
rect 146574 199552 146576 199572
rect 146576 199552 146628 199572
rect 146628 199552 146630 199572
rect 147034 199688 147090 199744
rect 148184 199858 148240 199914
rect 146666 193704 146722 193760
rect 146298 147736 146354 147792
rect 146942 196560 146998 196616
rect 146758 142704 146814 142760
rect 147310 199552 147366 199608
rect 147310 198464 147366 198520
rect 147402 198328 147458 198384
rect 147126 194248 147182 194304
rect 147862 199588 147864 199608
rect 147864 199588 147916 199608
rect 147916 199588 147918 199608
rect 147862 199552 147918 199588
rect 147586 192888 147642 192944
rect 147494 192752 147550 192808
rect 147310 189080 147366 189136
rect 147218 187176 147274 187232
rect 149012 199824 149068 199880
rect 148736 199688 148792 199744
rect 148230 196424 148286 196480
rect 148138 190984 148194 191040
rect 147310 139984 147366 140040
rect 148138 148280 148194 148336
rect 148690 197920 148746 197976
rect 148414 142840 148470 142896
rect 149058 199688 149114 199744
rect 149472 199824 149528 199880
rect 148966 197920 149022 197976
rect 149150 196696 149206 196752
rect 150300 199824 150356 199880
rect 149518 144064 149574 144120
rect 149702 182008 149758 182064
rect 149702 144200 149758 144256
rect 150254 199572 150310 199608
rect 150254 199552 150256 199572
rect 150256 199552 150308 199572
rect 150308 199552 150310 199572
rect 150254 199180 150256 199200
rect 150256 199180 150308 199200
rect 150308 199180 150310 199200
rect 150254 199144 150310 199180
rect 150668 199858 150724 199914
rect 150530 197376 150586 197432
rect 150438 191528 150494 191584
rect 150714 199572 150770 199608
rect 150714 199552 150716 199572
rect 150716 199552 150768 199572
rect 150768 199552 150770 199572
rect 150714 199008 150770 199064
rect 150990 199008 151046 199064
rect 150990 198464 151046 198520
rect 151082 198056 151138 198112
rect 151082 196696 151138 196752
rect 150898 189080 150954 189136
rect 151496 199688 151552 199744
rect 151956 199858 152012 199914
rect 152140 199858 152196 199914
rect 152324 199858 152380 199914
rect 152692 199824 152748 199880
rect 151910 199688 151966 199744
rect 152094 199688 152150 199744
rect 151450 199552 151506 199608
rect 151634 199552 151690 199608
rect 151634 199008 151690 199064
rect 151634 198872 151690 198928
rect 152094 199008 152150 199064
rect 151818 198872 151874 198928
rect 151726 197648 151782 197704
rect 151174 187312 151230 187368
rect 150070 145560 150126 145616
rect 152370 199688 152426 199744
rect 152646 199688 152702 199744
rect 152968 199858 153024 199914
rect 152278 198872 152334 198928
rect 152278 193976 152334 194032
rect 152462 189624 152518 189680
rect 152646 199144 152702 199200
rect 152738 198872 152794 198928
rect 152922 199552 152978 199608
rect 152646 196016 152702 196072
rect 152646 194520 152702 194576
rect 152646 189760 152702 189816
rect 153612 199858 153668 199914
rect 153382 199552 153438 199608
rect 153106 199180 153108 199200
rect 153108 199180 153160 199200
rect 153160 199180 153162 199200
rect 153106 199144 153162 199180
rect 153290 196424 153346 196480
rect 153290 196152 153346 196208
rect 153382 196016 153438 196072
rect 152554 148280 152610 148336
rect 153934 199688 153990 199744
rect 154532 199824 154588 199880
rect 153750 198872 153806 198928
rect 153934 199144 153990 199200
rect 153658 189624 153714 189680
rect 153566 188944 153622 189000
rect 153566 188536 153622 188592
rect 153474 186904 153530 186960
rect 153842 195472 153898 195528
rect 154118 193704 154174 193760
rect 154394 199588 154396 199608
rect 154396 199588 154448 199608
rect 154448 199588 154450 199608
rect 154394 199552 154450 199588
rect 154486 196016 154542 196072
rect 154394 139984 154450 140040
rect 155820 199858 155876 199914
rect 155774 199688 155830 199744
rect 156556 199858 156612 199914
rect 157016 199824 157072 199880
rect 157200 199858 157256 199914
rect 155866 191120 155922 191176
rect 156234 196424 156290 196480
rect 156602 199688 156658 199744
rect 156786 199724 156788 199744
rect 156788 199724 156840 199744
rect 156840 199724 156842 199744
rect 156786 199688 156842 199724
rect 156510 196696 156566 196752
rect 156418 196016 156474 196072
rect 157154 199552 157210 199608
rect 157890 199688 157946 199744
rect 158304 199858 158360 199914
rect 157890 198736 157946 198792
rect 158534 199688 158590 199744
rect 158258 199552 158314 199608
rect 158166 198872 158222 198928
rect 158948 199858 159004 199914
rect 158718 198056 158774 198112
rect 157982 144064 158038 144120
rect 157246 142296 157302 142352
rect 159224 199858 159280 199914
rect 159454 199688 159510 199744
rect 159960 199824 160016 199880
rect 159270 199552 159326 199608
rect 159270 197376 159326 197432
rect 159270 196968 159326 197024
rect 158902 182960 158958 183016
rect 159730 198500 159732 198520
rect 159732 198500 159784 198520
rect 159784 198500 159786 198520
rect 159730 198464 159786 198500
rect 159822 198192 159878 198248
rect 160236 199858 160292 199914
rect 160604 199858 160660 199914
rect 161248 199858 161304 199914
rect 160558 199688 160614 199744
rect 160742 199552 160798 199608
rect 160926 198328 160982 198384
rect 160834 197784 160890 197840
rect 161202 196696 161258 196752
rect 161478 199688 161534 199744
rect 161662 199688 161718 199744
rect 161938 198600 161994 198656
rect 162030 197376 162086 197432
rect 162628 199824 162684 199880
rect 162490 199280 162546 199336
rect 163548 199824 163604 199880
rect 163226 197920 163282 197976
rect 163226 197784 163282 197840
rect 163502 196968 163558 197024
rect 164008 199824 164064 199880
rect 163686 196696 163742 196752
rect 163594 189080 163650 189136
rect 164054 198908 164056 198928
rect 164056 198908 164108 198928
rect 164108 198908 164110 198928
rect 164054 198872 164110 198908
rect 164330 198464 164386 198520
rect 164238 197920 164294 197976
rect 164238 196560 164294 196616
rect 165204 199858 165260 199914
rect 164514 199552 164570 199608
rect 164882 199552 164938 199608
rect 164882 198872 164938 198928
rect 164790 198600 164846 198656
rect 165158 199688 165214 199744
rect 165664 199824 165720 199880
rect 164698 196696 164754 196752
rect 164514 195336 164570 195392
rect 165158 198736 165214 198792
rect 162766 140120 162822 140176
rect 164422 145560 164478 145616
rect 165434 198756 165490 198792
rect 165434 198736 165436 198756
rect 165436 198736 165488 198756
rect 165488 198736 165490 198756
rect 165434 197920 165490 197976
rect 165434 195200 165490 195256
rect 166032 199824 166088 199880
rect 166216 199824 166272 199880
rect 165894 199280 165950 199336
rect 165894 197376 165950 197432
rect 166584 199824 166640 199880
rect 166860 199858 166916 199914
rect 166814 199688 166870 199744
rect 167320 199858 167376 199914
rect 167504 199858 167560 199914
rect 167458 199688 167514 199744
rect 167090 198328 167146 198384
rect 167642 198872 167698 198928
rect 167642 197648 167698 197704
rect 168608 199824 168664 199880
rect 168102 197648 168158 197704
rect 168102 196288 168158 196344
rect 168010 193840 168066 193896
rect 168378 198872 168434 198928
rect 168654 199552 168710 199608
rect 169252 199824 169308 199880
rect 169436 199824 169492 199880
rect 169896 199858 169952 199914
rect 169390 199572 169446 199608
rect 169390 199552 169392 199572
rect 169392 199552 169444 199572
rect 169444 199552 169446 199572
rect 168838 191664 168894 191720
rect 168746 185952 168802 186008
rect 169850 199688 169906 199744
rect 170632 199858 170688 199914
rect 169666 196424 169722 196480
rect 168470 148416 168526 148472
rect 170310 199552 170366 199608
rect 170218 194928 170274 194984
rect 170908 199858 170964 199914
rect 170034 187584 170090 187640
rect 165618 141752 165674 141808
rect 169022 145696 169078 145752
rect 169758 143520 169814 143576
rect 141606 139304 141662 139360
rect 146666 139304 146722 139360
rect 154026 139304 154082 139360
rect 170862 199552 170918 199608
rect 170954 199280 171010 199336
rect 170954 198736 171010 198792
rect 170862 197512 170918 197568
rect 170770 197376 170826 197432
rect 170770 196852 170826 196888
rect 170770 196832 170772 196852
rect 170772 196832 170824 196852
rect 170824 196832 170826 196852
rect 170862 196696 170918 196752
rect 171322 199688 171378 199744
rect 171644 199858 171700 199914
rect 170954 195608 171010 195664
rect 172012 199858 172068 199914
rect 171690 199552 171746 199608
rect 171414 194792 171470 194848
rect 171690 199008 171746 199064
rect 172472 199858 172528 199914
rect 172748 199824 172804 199880
rect 173116 199824 173172 199880
rect 172334 198872 172390 198928
rect 172610 199416 172666 199472
rect 171506 145832 171562 145888
rect 172518 193160 172574 193216
rect 173070 196696 173126 196752
rect 172978 196424 173034 196480
rect 173852 199858 173908 199914
rect 173254 198600 173310 198656
rect 173346 196968 173402 197024
rect 173438 195744 173494 195800
rect 173852 199708 173908 199744
rect 174312 199858 174368 199914
rect 174496 199858 174552 199914
rect 174680 199858 174736 199914
rect 173852 199688 173854 199708
rect 173854 199688 173906 199708
rect 173906 199688 173908 199708
rect 173714 198600 173770 198656
rect 173714 193160 173770 193216
rect 173714 190712 173770 190768
rect 174542 199688 174598 199744
rect 174634 198600 174690 198656
rect 174542 196016 174598 196072
rect 174726 195744 174782 195800
rect 174726 192616 174782 192672
rect 175784 199858 175840 199914
rect 175738 197376 175794 197432
rect 175462 189080 175518 189136
rect 175646 186088 175702 186144
rect 176612 199858 176668 199914
rect 176888 199858 176944 199914
rect 176198 199416 176254 199472
rect 176382 193160 176438 193216
rect 176566 178608 176622 178664
rect 176566 146920 176622 146976
rect 178130 199960 178186 200016
rect 177394 196968 177450 197024
rect 177854 199824 177910 199880
rect 177670 198736 177726 198792
rect 178038 141616 178094 141672
rect 178590 199688 178646 199744
rect 178774 200368 178830 200424
rect 180430 200232 180486 200288
rect 180062 199960 180118 200016
rect 178866 199552 178922 199608
rect 178682 198872 178738 198928
rect 178590 194112 178646 194168
rect 178590 143384 178646 143440
rect 179326 199416 179382 199472
rect 179602 199008 179658 199064
rect 179418 197920 179474 197976
rect 179326 190984 179382 191040
rect 178866 142840 178922 142896
rect 179234 140256 179290 140312
rect 179418 142976 179474 143032
rect 179510 141480 179566 141536
rect 180522 200096 180578 200152
rect 180246 199688 180302 199744
rect 180062 198464 180118 198520
rect 179602 141344 179658 141400
rect 180706 199416 180762 199472
rect 180706 199008 180762 199064
rect 180246 198328 180302 198384
rect 183558 197920 183614 197976
rect 181810 195064 181866 195120
rect 182086 191392 182142 191448
rect 182086 191120 182142 191176
rect 181994 141888 182050 141944
rect 181902 141616 181958 141672
rect 182270 145968 182326 146024
rect 183374 184456 183430 184512
rect 184754 144336 184810 144392
rect 183466 142704 183522 142760
rect 183374 141480 183430 141536
rect 183282 140528 183338 140584
rect 184662 142568 184718 142624
rect 184846 140664 184902 140720
rect 186226 143112 186282 143168
rect 186134 140392 186190 140448
rect 182178 139440 182234 139496
rect 186318 139440 186374 139496
rect 187146 191120 187202 191176
rect 187146 190848 187202 190904
rect 186778 143384 186834 143440
rect 186962 143384 187018 143440
rect 186594 142976 186650 143032
rect 186778 142976 186834 143032
rect 186594 142432 186650 142488
rect 187146 139712 187202 139768
rect 187514 144200 187570 144256
rect 187422 139576 187478 139632
rect 187606 143112 187662 143168
rect 187514 139440 187570 139496
rect 180522 139304 180578 139360
rect 180706 139304 180762 139360
rect 186410 139304 186466 139360
rect 187054 139304 187110 139360
rect 123482 80552 123538 80608
rect 122286 78512 122342 78568
rect 124586 78376 124642 78432
rect 123482 71712 123538 71768
rect 131854 80316 131856 80336
rect 131856 80316 131908 80336
rect 131908 80316 131910 80336
rect 127438 79736 127494 79792
rect 131854 80280 131910 80316
rect 128450 78512 128506 78568
rect 132222 80180 132224 80200
rect 132224 80180 132276 80200
rect 132276 80180 132278 80200
rect 132222 80144 132278 80180
rect 131854 80008 131910 80064
rect 129002 79636 129004 79656
rect 129004 79636 129056 79656
rect 129056 79636 129058 79656
rect 129002 79600 129058 79636
rect 128634 78240 128690 78296
rect 128450 74432 128506 74488
rect 131026 72664 131082 72720
rect 132636 79906 132692 79962
rect 132498 79600 132554 79656
rect 132820 79736 132876 79792
rect 133188 79906 133244 79962
rect 132590 75928 132646 75984
rect 132866 79600 132922 79656
rect 132682 67224 132738 67280
rect 134016 79872 134072 79928
rect 134384 79872 134440 79928
rect 133510 74160 133566 74216
rect 134338 79736 134394 79792
rect 134660 79906 134716 79962
rect 134660 79772 134662 79792
rect 134662 79772 134714 79792
rect 134714 79772 134716 79792
rect 134660 79736 134716 79772
rect 135120 79872 135176 79928
rect 134936 79736 134992 79792
rect 135856 79872 135912 79928
rect 135304 79736 135360 79792
rect 136408 79906 136464 79962
rect 136684 79906 136740 79962
rect 134614 78512 134670 78568
rect 134614 78104 134670 78160
rect 134890 77968 134946 78024
rect 135074 78376 135130 78432
rect 135902 79772 135904 79792
rect 135904 79772 135956 79792
rect 135956 79772 135958 79792
rect 135902 79736 135958 79772
rect 135626 79056 135682 79112
rect 135718 77152 135774 77208
rect 134798 64504 134854 64560
rect 134798 63824 134854 63880
rect 136592 79770 136648 79826
rect 136960 79906 137016 79962
rect 137328 79906 137384 79962
rect 137512 79906 137568 79962
rect 137696 79906 137752 79962
rect 138248 79906 138304 79962
rect 138432 79906 138488 79962
rect 137972 79838 138028 79894
rect 138616 79906 138672 79962
rect 136638 79056 136694 79112
rect 136638 76744 136694 76800
rect 136086 76064 136142 76120
rect 135902 70216 135958 70272
rect 135810 68856 135866 68912
rect 136362 75928 136418 75984
rect 136730 75112 136786 75168
rect 137190 79600 137246 79656
rect 137098 77696 137154 77752
rect 136914 66136 136970 66192
rect 137650 79736 137706 79792
rect 137374 79192 137430 79248
rect 137466 78920 137522 78976
rect 137742 79600 137798 79656
rect 137742 77560 137798 77616
rect 138294 79736 138350 79792
rect 139260 79872 139316 79928
rect 139444 79872 139500 79928
rect 139168 79736 139224 79792
rect 139306 79736 139362 79792
rect 139720 79906 139776 79962
rect 138478 79600 138534 79656
rect 138386 79328 138442 79384
rect 138662 79600 138718 79656
rect 138754 77560 138810 77616
rect 138662 76880 138718 76936
rect 139122 79328 139178 79384
rect 139306 79192 139362 79248
rect 138846 67496 138902 67552
rect 140088 79872 140144 79928
rect 139950 79736 140006 79792
rect 140272 79906 140328 79962
rect 139398 74432 139454 74488
rect 139582 76336 139638 76392
rect 140640 79872 140696 79928
rect 140916 79872 140972 79928
rect 140134 79328 140190 79384
rect 140042 77832 140098 77888
rect 140778 79484 140834 79520
rect 140778 79464 140780 79484
rect 140780 79464 140832 79484
rect 140832 79464 140834 79484
rect 140686 79328 140742 79384
rect 140226 76744 140282 76800
rect 139766 66952 139822 67008
rect 140778 79192 140834 79248
rect 141422 79636 141424 79656
rect 141424 79636 141476 79656
rect 141476 79636 141478 79656
rect 141238 79464 141294 79520
rect 141238 79192 141294 79248
rect 141238 78104 141294 78160
rect 141422 79600 141478 79636
rect 141698 69944 141754 70000
rect 141606 68720 141662 68776
rect 141514 68584 141570 68640
rect 140962 66000 141018 66056
rect 140870 65728 140926 65784
rect 142940 79872 142996 79928
rect 142342 79056 142398 79112
rect 142066 70352 142122 70408
rect 142066 68312 142122 68368
rect 142802 79056 142858 79112
rect 143078 78376 143134 78432
rect 143492 79906 143548 79962
rect 143492 79736 143548 79792
rect 143722 79736 143778 79792
rect 143446 78512 143502 78568
rect 143814 72528 143870 72584
rect 144274 79736 144330 79792
rect 144366 78784 144422 78840
rect 144366 78104 144422 78160
rect 144780 79872 144836 79928
rect 145240 79906 145296 79962
rect 144826 79600 144882 79656
rect 144458 77832 144514 77888
rect 144826 79464 144882 79520
rect 145102 79600 145158 79656
rect 145010 78376 145066 78432
rect 144550 76472 144606 76528
rect 145286 79600 145342 79656
rect 145194 74976 145250 75032
rect 145608 79906 145664 79962
rect 145884 79906 145940 79962
rect 146160 79906 146216 79962
rect 146344 79838 146400 79894
rect 145562 79620 145618 79656
rect 145562 79600 145564 79620
rect 145564 79600 145616 79620
rect 145616 79600 145618 79620
rect 145470 79328 145526 79384
rect 145654 75792 145710 75848
rect 146022 77968 146078 78024
rect 146298 79600 146354 79656
rect 145562 72392 145618 72448
rect 147080 79872 147136 79928
rect 146758 79464 146814 79520
rect 147448 79906 147504 79962
rect 147632 79906 147688 79962
rect 146942 73752 146998 73808
rect 147586 79736 147642 79792
rect 147310 77968 147366 78024
rect 147034 71440 147090 71496
rect 148552 79872 148608 79928
rect 148276 79770 148332 79826
rect 149104 79872 149160 79928
rect 149472 79906 149528 79962
rect 149748 79906 149804 79962
rect 150024 79872 150080 79928
rect 149978 79736 150034 79792
rect 150208 79838 150264 79894
rect 150392 79838 150448 79894
rect 150668 79872 150724 79928
rect 148046 79600 148102 79656
rect 148230 79636 148232 79656
rect 148232 79636 148284 79656
rect 148284 79636 148286 79656
rect 148230 79600 148286 79636
rect 147954 76608 148010 76664
rect 148414 79464 148470 79520
rect 148598 78240 148654 78296
rect 148414 75520 148470 75576
rect 148966 79600 149022 79656
rect 149150 79600 149206 79656
rect 149518 79328 149574 79384
rect 149426 77968 149482 78024
rect 150346 79600 150402 79656
rect 150254 77968 150310 78024
rect 151220 79872 151276 79928
rect 151496 79906 151552 79962
rect 150622 78104 150678 78160
rect 150438 72936 150494 72992
rect 151174 78240 151230 78296
rect 150898 74024 150954 74080
rect 150622 69400 150678 69456
rect 151864 79906 151920 79962
rect 152140 79906 152196 79962
rect 152324 79906 152380 79962
rect 152600 79872 152656 79928
rect 153060 79872 153116 79928
rect 153336 79906 153392 79962
rect 153520 79906 153576 79962
rect 151358 79464 151414 79520
rect 151634 79600 151690 79656
rect 151542 77560 151598 77616
rect 152370 79736 152426 79792
rect 152508 79736 152564 79792
rect 151910 79600 151966 79656
rect 151726 77696 151782 77752
rect 151174 64640 151230 64696
rect 152278 79600 152334 79656
rect 153704 79906 153760 79962
rect 153888 79906 153944 79962
rect 154072 79872 154128 79928
rect 152554 79600 152610 79656
rect 152462 71712 152518 71768
rect 152186 70080 152242 70136
rect 152646 71712 152702 71768
rect 153290 77968 153346 78024
rect 153106 73616 153162 73672
rect 154440 79906 154496 79962
rect 154716 79906 154772 79962
rect 155176 79906 155232 79962
rect 155544 79906 155600 79962
rect 154026 79600 154082 79656
rect 153750 78920 153806 78976
rect 153566 74976 153622 75032
rect 153474 69400 153530 69456
rect 154762 79636 154764 79656
rect 154764 79636 154816 79656
rect 154816 79636 154818 79656
rect 154762 79600 154818 79636
rect 154762 79464 154818 79520
rect 154670 77152 154726 77208
rect 155406 76336 155462 76392
rect 156418 78648 156474 78704
rect 156602 78512 156658 78568
rect 156602 73072 156658 73128
rect 156510 71712 156566 71768
rect 156510 71032 156566 71088
rect 156878 79056 156934 79112
rect 156694 71712 156750 71768
rect 157154 79600 157210 79656
rect 157568 79872 157624 79928
rect 157844 79906 157900 79962
rect 157430 66680 157486 66736
rect 157890 79736 157946 79792
rect 158212 79906 158268 79962
rect 157982 78240 158038 78296
rect 158166 79772 158168 79792
rect 158168 79772 158220 79792
rect 158220 79772 158222 79792
rect 158166 79736 158222 79772
rect 158856 79736 158912 79792
rect 158074 76608 158130 76664
rect 159270 79736 159326 79792
rect 158442 76608 158498 76664
rect 158810 75928 158866 75984
rect 159270 79600 159326 79656
rect 159638 79328 159694 79384
rect 159822 77016 159878 77072
rect 160972 79872 161028 79928
rect 161156 79872 161212 79928
rect 160098 75792 160154 75848
rect 160006 73752 160062 73808
rect 159730 71576 159786 71632
rect 159362 68856 159418 68912
rect 158994 65456 159050 65512
rect 158810 64776 158866 64832
rect 160374 79464 160430 79520
rect 162076 79906 162132 79962
rect 160466 75928 160522 75984
rect 161110 78648 161166 78704
rect 161524 79736 161580 79792
rect 161938 79736 161994 79792
rect 161478 79600 161534 79656
rect 162904 79906 162960 79962
rect 162030 77152 162086 77208
rect 162582 79464 162638 79520
rect 162950 79600 163006 79656
rect 162674 78512 162730 78568
rect 163456 79906 163512 79962
rect 163916 79872 163972 79928
rect 164284 79872 164340 79928
rect 164468 79872 164524 79928
rect 163134 67496 163190 67552
rect 165112 79906 165168 79962
rect 165296 79906 165352 79962
rect 165480 79872 165536 79928
rect 165848 79906 165904 79962
rect 166032 79906 166088 79962
rect 163870 78376 163926 78432
rect 164146 79600 164202 79656
rect 164606 78512 164662 78568
rect 165250 79736 165306 79792
rect 165066 79600 165122 79656
rect 164974 76608 165030 76664
rect 164882 76472 164938 76528
rect 165710 79736 165766 79792
rect 165618 79600 165674 79656
rect 165250 72800 165306 72856
rect 165986 79736 166042 79792
rect 165802 77968 165858 78024
rect 165342 68312 165398 68368
rect 166584 79906 166640 79962
rect 167044 79906 167100 79962
rect 167412 79872 167468 79928
rect 167872 79872 167928 79928
rect 165986 78512 166042 78568
rect 166538 79620 166594 79656
rect 166538 79600 166540 79620
rect 166540 79600 166592 79620
rect 166592 79600 166594 79620
rect 166170 71032 166226 71088
rect 166952 79736 167008 79792
rect 168056 79736 168112 79792
rect 168240 79872 168296 79928
rect 168608 79906 168664 79962
rect 167826 78920 167882 78976
rect 168378 79192 168434 79248
rect 168286 78920 168342 78976
rect 168746 79600 168802 79656
rect 168654 68584 168710 68640
rect 169252 79906 169308 79962
rect 169620 79872 169676 79928
rect 169482 78784 169538 78840
rect 169988 79906 170044 79962
rect 170264 79906 170320 79962
rect 170724 79872 170780 79928
rect 169758 76064 169814 76120
rect 170034 75928 170090 75984
rect 169666 72392 169722 72448
rect 171092 79872 171148 79928
rect 170862 78920 170918 78976
rect 171138 79736 171194 79792
rect 171230 79600 171286 79656
rect 171230 79192 171286 79248
rect 171598 79736 171654 79792
rect 171920 79838 171976 79894
rect 172288 79906 172344 79962
rect 172472 79906 172528 79962
rect 172656 79872 172712 79928
rect 170954 73072 171010 73128
rect 171138 68720 171194 68776
rect 171966 75928 172022 75984
rect 171322 69672 171378 69728
rect 172518 79736 172574 79792
rect 173116 79906 173172 79962
rect 172702 78920 172758 78976
rect 173070 79736 173126 79792
rect 173070 78104 173126 78160
rect 173162 75520 173218 75576
rect 173070 71168 173126 71224
rect 172058 68348 172060 68368
rect 172060 68348 172112 68368
rect 172112 68348 172114 68368
rect 172058 68312 172114 68348
rect 173944 79906 174000 79962
rect 173806 75656 173862 75712
rect 173898 72936 173954 72992
rect 173530 68312 173586 68368
rect 174818 79736 174874 79792
rect 174726 79328 174782 79384
rect 174726 78140 174728 78160
rect 174728 78140 174780 78160
rect 174780 78140 174782 78160
rect 174726 78104 174782 78140
rect 174634 76472 174690 76528
rect 174634 67360 174690 67416
rect 175968 79906 176024 79962
rect 176336 79906 176392 79962
rect 175094 78376 175150 78432
rect 175370 79328 175426 79384
rect 176014 75792 176070 75848
rect 176750 79736 176806 79792
rect 176198 75248 176254 75304
rect 176474 68176 176530 68232
rect 177256 79736 177312 79792
rect 177302 76744 177358 76800
rect 177578 78512 177634 78568
rect 177946 80552 178002 80608
rect 179234 80416 179290 80472
rect 177946 79872 178002 79928
rect 177946 76472 178002 76528
rect 179602 80008 179658 80064
rect 186318 80552 186374 80608
rect 185582 80416 185638 80472
rect 179050 77696 179106 77752
rect 179970 77832 180026 77888
rect 178958 75384 179014 75440
rect 186318 79056 186374 79112
rect 183926 78376 183982 78432
rect 184202 78376 184258 78432
rect 186318 78376 186374 78432
rect 182178 78104 182234 78160
rect 181442 74296 181498 74352
rect 186962 70216 187018 70272
rect 188434 80416 188490 80472
rect 188618 80144 188674 80200
rect 189078 195200 189134 195256
rect 189078 194792 189134 194848
rect 188894 139984 188950 140040
rect 188986 91160 189042 91216
rect 188434 74432 188490 74488
rect 188986 66136 189042 66192
rect 189722 199552 189778 199608
rect 189998 197512 190054 197568
rect 189906 195200 189962 195256
rect 190458 142296 190514 142352
rect 189906 136584 189962 136640
rect 189998 81368 190054 81424
rect 189998 80416 190054 80472
rect 189630 77152 189686 77208
rect 191194 200640 191250 200696
rect 191194 82728 191250 82784
rect 192114 142976 192170 143032
rect 192206 139304 192262 139360
rect 192390 143520 192446 143576
rect 192666 141888 192722 141944
rect 192574 140392 192630 140448
rect 192850 143520 192906 143576
rect 192574 72664 192630 72720
rect 192206 66952 192262 67008
rect 193586 142432 193642 142488
rect 194598 195336 194654 195392
rect 193954 80824 194010 80880
rect 195426 259528 195482 259584
rect 195334 145832 195390 145888
rect 196622 263608 196678 263664
rect 195426 142568 195482 142624
rect 195242 139168 195298 139224
rect 195426 137400 195482 137456
rect 195426 78240 195482 78296
rect 196990 145560 197046 145616
rect 197358 197920 197414 197976
rect 197910 140664 197966 140720
rect 197726 139032 197782 139088
rect 198830 196424 198886 196480
rect 198830 192888 198886 192944
rect 198830 72528 198886 72584
rect 199198 74976 199254 75032
rect 200118 187448 200174 187504
rect 199474 138624 199530 138680
rect 199382 81232 199438 81288
rect 202234 194112 202290 194168
rect 201590 192752 201646 192808
rect 200394 76472 200450 76528
rect 200578 73888 200634 73944
rect 200210 66972 200266 67008
rect 200210 66952 200212 66972
rect 200212 66952 200264 66972
rect 200264 66952 200266 66972
rect 200762 137264 200818 137320
rect 199474 65592 199530 65648
rect 201038 191256 201094 191312
rect 200854 134408 200910 134464
rect 200946 81776 201002 81832
rect 201038 67224 201094 67280
rect 200762 64640 200818 64696
rect 201498 187040 201554 187096
rect 201498 71440 201554 71496
rect 201498 70216 201554 70272
rect 201590 67088 201646 67144
rect 202878 81096 202934 81152
rect 203522 148416 203578 148472
rect 203430 80960 203486 81016
rect 204258 70216 204314 70272
rect 204350 69944 204406 70000
rect 204626 68312 204682 68368
rect 205086 81640 205142 81696
rect 205638 69944 205694 70000
rect 205822 68856 205878 68912
rect 206098 68176 206154 68232
rect 207110 71440 207166 71496
rect 207478 187176 207534 187232
rect 207478 81232 207534 81288
rect 207754 141752 207810 141808
rect 208674 185680 208730 185736
rect 209042 188536 209098 188592
rect 209042 75792 209098 75848
rect 211158 194928 211214 194984
rect 209962 76764 210018 76800
rect 209962 76744 209964 76764
rect 209964 76744 210016 76764
rect 210016 76744 210018 76764
rect 209870 68720 209926 68776
rect 210330 75248 210386 75304
rect 211158 66816 211214 66872
rect 212446 195744 212502 195800
rect 211526 195608 211582 195664
rect 212446 194928 212502 194984
rect 211434 77696 211490 77752
rect 211342 63416 211398 63472
rect 211250 63144 211306 63200
rect 212814 79328 212870 79384
rect 212630 75520 212686 75576
rect 213090 78512 213146 78568
rect 214102 192616 214158 192672
rect 214010 75656 214066 75712
rect 214194 178880 214250 178936
rect 214378 189760 214434 189816
rect 214562 187448 214618 187504
rect 214562 186768 214618 186824
rect 214378 78920 214434 78976
rect 214470 78784 214526 78840
rect 214194 63280 214250 63336
rect 215390 76336 215446 76392
rect 218058 195472 218114 195528
rect 214838 65320 214894 65376
rect 215942 77832 215998 77888
rect 215758 65864 215814 65920
rect 216126 148280 216182 148336
rect 217046 185816 217102 185872
rect 216862 181328 216918 181384
rect 216770 81912 216826 81968
rect 217322 184320 217378 184376
rect 217230 183368 217286 183424
rect 217414 80688 217470 80744
rect 217322 78648 217378 78704
rect 217230 77016 217286 77072
rect 217046 72936 217102 72992
rect 216954 69536 217010 69592
rect 218518 188264 218574 188320
rect 218150 183232 218206 183288
rect 218242 183096 218298 183152
rect 218242 182552 218298 182608
rect 218242 70896 218298 70952
rect 218518 76880 218574 76936
rect 218150 66000 218206 66056
rect 216862 65728 216918 65784
rect 220082 195608 220138 195664
rect 224222 192752 224278 192808
rect 237378 193976 237434 194032
rect 242162 188944 242218 189000
rect 263598 268368 263654 268424
rect 282918 186224 282974 186280
rect 309138 182688 309194 182744
rect 340878 194248 340934 194304
rect 374642 201048 374698 201104
rect 371238 189896 371294 189952
rect 378138 188400 378194 188456
rect 386418 195744 386474 195800
rect 420918 196832 420974 196888
rect 425058 194384 425114 194440
rect 416778 191528 416834 191584
rect 440238 191392 440294 191448
rect 445022 197104 445078 197160
rect 444378 184456 444434 184512
rect 409878 183504 409934 183560
rect 466458 201728 466514 201784
rect 463698 183368 463754 183424
rect 459558 182008 459614 182064
rect 485778 195880 485834 195936
rect 489918 183232 489974 183288
rect 509238 200912 509294 200968
rect 520278 262656 520334 262712
rect 516138 191256 516194 191312
rect 535458 269728 535514 269784
rect 542358 194520 542414 194576
rect 539598 181328 539654 181384
rect 494702 180376 494758 180432
rect 481638 180240 481694 180296
rect 546498 188264 546554 188320
rect 544474 177928 544530 177984
rect 548614 199552 548670 199608
rect 552662 184184 552718 184240
rect 548522 176568 548578 176624
rect 556894 178608 556950 178664
rect 558918 195064 558974 195120
rect 561034 184320 561090 184376
rect 561678 200776 561734 200832
rect 565082 182960 565138 183016
rect 566554 189760 566610 189816
rect 566646 187448 566702 187504
rect 566462 187312 566518 187368
rect 567842 191120 567898 191176
rect 569314 186904 569370 186960
rect 567934 185816 567990 185872
rect 565174 180512 565230 180568
rect 571982 195336 572038 195392
rect 572166 187176 572222 187232
rect 570786 185680 570842 185736
rect 570694 178880 570750 178936
rect 574834 192616 574890 192672
rect 574926 190304 574982 190360
rect 580170 702500 580226 702536
rect 580170 702480 580172 702500
rect 580172 702480 580224 702500
rect 580224 702480 580226 702500
rect 580170 698400 580226 698456
rect 580170 694320 580226 694376
rect 579802 686160 579858 686216
rect 576122 196696 576178 196752
rect 576306 196560 576362 196616
rect 577502 195200 577558 195256
rect 576214 190984 576270 191040
rect 575110 189624 575166 189680
rect 575018 187040 575074 187096
rect 573362 178744 573418 178800
rect 580170 678000 580226 678056
rect 580170 669840 580226 669896
rect 580170 665760 580226 665816
rect 579986 649440 580042 649496
rect 580170 645360 580226 645416
rect 580170 633800 580226 633856
rect 580170 629720 580226 629776
rect 580538 625640 580594 625696
rect 580170 609320 580226 609376
rect 580354 605240 580410 605296
rect 580170 597080 580226 597136
rect 580170 593000 580226 593056
rect 580170 584840 580226 584896
rect 578882 577360 578938 577416
rect 578238 192480 578294 192536
rect 580170 573280 580226 573336
rect 579710 569200 579766 569256
rect 580170 565120 580226 565176
rect 579618 561040 579674 561096
rect 580078 548800 580134 548856
rect 580170 544720 580226 544776
rect 579710 540640 579766 540696
rect 580170 536560 580226 536616
rect 580170 528400 580226 528456
rect 580170 524320 580226 524376
rect 579710 520920 579766 520976
rect 580170 516840 580226 516896
rect 579618 512760 579674 512816
rect 580170 508680 580226 508736
rect 580078 504600 580134 504656
rect 580170 500520 580226 500576
rect 580170 496440 580226 496496
rect 580170 488280 580226 488336
rect 580170 484200 580226 484256
rect 580170 480120 580226 480176
rect 580170 476040 580226 476096
rect 580170 471996 580172 472016
rect 580172 471996 580224 472016
rect 580224 471996 580226 472016
rect 580170 471960 580226 471996
rect 580170 467900 580226 467936
rect 580170 467880 580172 467900
rect 580172 467880 580224 467900
rect 580224 467880 580226 467900
rect 580170 463800 580226 463856
rect 580170 460400 580226 460456
rect 580078 456320 580134 456376
rect 580170 452240 580226 452296
rect 579710 448160 579766 448216
rect 580170 444080 580226 444136
rect 580170 435920 580226 435976
rect 580170 431840 580226 431896
rect 580170 427760 580226 427816
rect 580170 423700 580226 423736
rect 580170 423680 580172 423700
rect 580172 423680 580224 423700
rect 580224 423680 580226 423700
rect 580170 419600 580226 419656
rect 580170 415520 580226 415576
rect 579986 411440 580042 411496
rect 580170 407360 580226 407416
rect 580170 403960 580226 404016
rect 579710 399880 579766 399936
rect 580170 395800 580226 395856
rect 580170 391720 580226 391776
rect 580170 387640 580226 387696
rect 578974 383560 579030 383616
rect 580170 375420 580226 375456
rect 580170 375400 580172 375420
rect 580172 375400 580224 375420
rect 580224 375400 580226 375420
rect 579802 371320 579858 371376
rect 580170 367240 580226 367296
rect 580170 359080 580226 359136
rect 580170 355000 580226 355056
rect 580170 350920 580226 350976
rect 580170 346840 580226 346896
rect 579710 343440 579766 343496
rect 579618 339360 579674 339416
rect 579710 331236 579712 331256
rect 579712 331236 579764 331256
rect 579764 331236 579766 331256
rect 579710 331200 579766 331236
rect 579066 323040 579122 323096
rect 579710 318960 579766 319016
rect 579618 314880 579674 314936
rect 580170 310800 580226 310856
rect 580170 306720 580226 306776
rect 580170 302640 580226 302696
rect 579158 298560 579214 298616
rect 580170 294480 580226 294536
rect 579986 290400 580042 290456
rect 579986 286320 580042 286376
rect 580170 282940 580226 282976
rect 580170 282920 580172 282940
rect 580172 282920 580224 282940
rect 580224 282920 580226 282940
rect 580170 278840 580226 278896
rect 580170 274760 580226 274816
rect 579710 270680 579766 270736
rect 579618 266600 579674 266656
rect 580262 262520 580318 262576
rect 580262 258440 580318 258496
rect 579802 254360 579858 254416
rect 579986 250280 580042 250336
rect 580170 242120 580226 242176
rect 580170 238040 580226 238096
rect 579986 225800 580042 225856
rect 580170 197920 580226 197976
rect 580538 588920 580594 588976
rect 580446 379480 580502 379536
rect 580354 199280 580410 199336
rect 580262 197240 580318 197296
rect 579802 193840 579858 193896
rect 579618 189760 579674 189816
rect 580262 185680 580318 185736
rect 580170 181600 580226 181656
rect 580170 177520 580226 177576
rect 558274 176432 558330 176488
rect 544382 176296 544438 176352
rect 382278 176160 382334 176216
rect 367098 176024 367154 176080
rect 351918 175888 351974 175944
rect 580170 173440 580226 173496
rect 580262 169360 580318 169416
rect 580170 165280 580226 165336
rect 580170 161880 580226 161936
rect 579618 153720 579674 153776
rect 580170 149676 580172 149696
rect 580172 149676 580224 149696
rect 580224 149676 580226 149696
rect 580170 149640 580226 149676
rect 580170 145560 580226 145616
rect 579618 142704 579674 142760
rect 580170 137400 580226 137456
rect 580170 125160 580226 125216
rect 580170 112920 580226 112976
rect 580170 85040 580226 85096
rect 580630 327120 580686 327176
rect 580538 199416 580594 199472
rect 580722 229880 580778 229936
rect 580814 214240 580870 214296
rect 580906 210160 580962 210216
rect 582378 690240 582434 690296
rect 581734 661680 581790 661736
rect 581642 657600 581698 657656
rect 580998 185544 581054 185600
rect 581826 440000 581882 440056
rect 581734 193976 581790 194032
rect 582470 682080 582526 682136
rect 582654 637880 582710 637936
rect 582562 621560 582618 621616
rect 582838 617480 582894 617536
rect 582746 613400 582802 613456
rect 582654 200640 582710 200696
rect 582930 556960 582986 557016
rect 582838 195472 582894 195528
rect 582562 183096 582618 183152
rect 582470 182824 582526 182880
rect 583022 532480 583078 532536
rect 582930 180648 582986 180704
rect 580538 147736 580594 147792
rect 580446 141480 580502 141536
rect 580354 129240 580410 129296
rect 580722 133320 580778 133376
rect 580630 121080 580686 121136
rect 580538 117000 580594 117056
rect 580446 108840 580502 108896
rect 580354 104760 580410 104816
rect 580262 72800 580318 72856
rect 579986 68720 580042 68776
rect 580630 101360 580686 101416
rect 580446 97280 580502 97336
rect 580538 89120 580594 89176
rect 580722 93200 580778 93256
rect 580630 76880 580686 76936
rect 580722 72256 580778 72312
rect 580446 62056 580502 62112
rect 580170 48320 580226 48376
rect 579986 44240 580042 44296
rect 580170 40840 580226 40896
rect 580170 36760 580226 36816
rect 580170 32680 580226 32736
rect 580170 24520 580226 24576
rect 580170 20440 580226 20496
rect 580170 16360 580226 16416
rect 580170 12280 580226 12336
rect 580170 8236 580172 8256
rect 580172 8236 580224 8256
rect 580224 8236 580226 8256
rect 580170 8200 580226 8236
rect 580170 4120 580226 4176
rect 578882 40 578938 96
<< metal3 >>
rect 580165 702538 580231 702541
rect 583520 702538 584960 702628
rect 580165 702536 584960 702538
rect 580165 702480 580170 702536
rect 580226 702480 584960 702536
rect 580165 702478 584960 702480
rect 580165 702475 580231 702478
rect 583520 702388 584960 702478
rect -960 701858 480 701948
rect 3049 701858 3115 701861
rect -960 701856 3115 701858
rect -960 701800 3054 701856
rect 3110 701800 3115 701856
rect -960 701798 3115 701800
rect -960 701708 480 701798
rect 3049 701795 3115 701798
rect 580165 698458 580231 698461
rect 583520 698458 584960 698548
rect 580165 698456 584960 698458
rect 580165 698400 580170 698456
rect 580226 698400 584960 698456
rect 580165 698398 584960 698400
rect 580165 698395 580231 698398
rect 583520 698308 584960 698398
rect -960 697628 480 697868
rect 580165 694378 580231 694381
rect 583520 694378 584960 694468
rect 580165 694376 584960 694378
rect 580165 694320 580170 694376
rect 580226 694320 584960 694376
rect 580165 694318 584960 694320
rect 580165 694315 580231 694318
rect 583520 694228 584960 694318
rect -960 693698 480 693788
rect 3141 693698 3207 693701
rect -960 693696 3207 693698
rect -960 693640 3146 693696
rect 3202 693640 3207 693696
rect -960 693638 3207 693640
rect -960 693548 480 693638
rect 3141 693635 3207 693638
rect 582373 690298 582439 690301
rect 583520 690298 584960 690388
rect 582373 690296 584960 690298
rect 582373 690240 582378 690296
rect 582434 690240 584960 690296
rect 582373 690238 584960 690240
rect 582373 690235 582439 690238
rect 583520 690148 584960 690238
rect -960 689618 480 689708
rect 3417 689618 3483 689621
rect -960 689616 3483 689618
rect -960 689560 3422 689616
rect 3478 689560 3483 689616
rect -960 689558 3483 689560
rect -960 689468 480 689558
rect 3417 689555 3483 689558
rect 579797 686218 579863 686221
rect 583520 686218 584960 686308
rect 579797 686216 584960 686218
rect 579797 686160 579802 686216
rect 579858 686160 584960 686216
rect 579797 686158 584960 686160
rect 579797 686155 579863 686158
rect 583520 686068 584960 686158
rect -960 685538 480 685628
rect 3141 685538 3207 685541
rect -960 685536 3207 685538
rect -960 685480 3146 685536
rect 3202 685480 3207 685536
rect -960 685478 3207 685480
rect -960 685388 480 685478
rect 3141 685475 3207 685478
rect 582465 682138 582531 682141
rect 583520 682138 584960 682228
rect 582465 682136 584960 682138
rect 582465 682080 582470 682136
rect 582526 682080 584960 682136
rect 582465 682078 584960 682080
rect 582465 682075 582531 682078
rect 583520 681988 584960 682078
rect -960 681458 480 681548
rect 3417 681458 3483 681461
rect -960 681456 3483 681458
rect -960 681400 3422 681456
rect 3478 681400 3483 681456
rect -960 681398 3483 681400
rect -960 681308 480 681398
rect 3417 681395 3483 681398
rect 580165 678058 580231 678061
rect 583520 678058 584960 678148
rect 580165 678056 584960 678058
rect 580165 678000 580170 678056
rect 580226 678000 584960 678056
rect 580165 677998 584960 678000
rect 580165 677995 580231 677998
rect 583520 677908 584960 677998
rect -960 677228 480 677468
rect 583520 673828 584960 674068
rect -960 673298 480 673388
rect 3233 673298 3299 673301
rect -960 673296 3299 673298
rect -960 673240 3238 673296
rect 3294 673240 3299 673296
rect -960 673238 3299 673240
rect -960 673148 480 673238
rect 3233 673235 3299 673238
rect 580165 669898 580231 669901
rect 583520 669898 584960 669988
rect 580165 669896 584960 669898
rect 580165 669840 580170 669896
rect 580226 669840 584960 669896
rect 580165 669838 584960 669840
rect 580165 669835 580231 669838
rect 583520 669748 584960 669838
rect -960 669218 480 669308
rect 3417 669218 3483 669221
rect -960 669216 3483 669218
rect -960 669160 3422 669216
rect 3478 669160 3483 669216
rect -960 669158 3483 669160
rect -960 669068 480 669158
rect 3417 669155 3483 669158
rect 580165 665818 580231 665821
rect 583520 665818 584960 665908
rect 580165 665816 584960 665818
rect 580165 665760 580170 665816
rect 580226 665760 584960 665816
rect 580165 665758 584960 665760
rect 580165 665755 580231 665758
rect 583520 665668 584960 665758
rect -960 665138 480 665228
rect 3233 665138 3299 665141
rect -960 665136 3299 665138
rect -960 665080 3238 665136
rect 3294 665080 3299 665136
rect -960 665078 3299 665080
rect -960 664988 480 665078
rect 3233 665075 3299 665078
rect 581729 661738 581795 661741
rect 583520 661738 584960 661828
rect 581729 661736 584960 661738
rect 581729 661680 581734 661736
rect 581790 661680 584960 661736
rect 581729 661678 584960 661680
rect 581729 661675 581795 661678
rect 583520 661588 584960 661678
rect -960 661058 480 661148
rect 3417 661058 3483 661061
rect -960 661056 3483 661058
rect -960 661000 3422 661056
rect 3478 661000 3483 661056
rect -960 660998 3483 661000
rect -960 660908 480 660998
rect 3417 660995 3483 660998
rect -960 657508 480 657748
rect 581637 657658 581703 657661
rect 583520 657658 584960 657748
rect 581637 657656 584960 657658
rect 581637 657600 581642 657656
rect 581698 657600 584960 657656
rect 581637 657598 584960 657600
rect 581637 657595 581703 657598
rect 583520 657508 584960 657598
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 583520 653428 584960 653668
rect -960 649348 480 649588
rect 579981 649498 580047 649501
rect 583520 649498 584960 649588
rect 579981 649496 584960 649498
rect 579981 649440 579986 649496
rect 580042 649440 584960 649496
rect 579981 649438 584960 649440
rect 579981 649435 580047 649438
rect 583520 649348 584960 649438
rect -960 645418 480 645508
rect 3417 645418 3483 645421
rect -960 645416 3483 645418
rect -960 645360 3422 645416
rect 3478 645360 3483 645416
rect -960 645358 3483 645360
rect -960 645268 480 645358
rect 3417 645355 3483 645358
rect 580165 645418 580231 645421
rect 583520 645418 584960 645508
rect 580165 645416 584960 645418
rect 580165 645360 580170 645416
rect 580226 645360 584960 645416
rect 580165 645358 584960 645360
rect 580165 645355 580231 645358
rect 583520 645268 584960 645358
rect 583520 641868 584960 642108
rect -960 641188 480 641428
rect 582649 637938 582715 637941
rect 583520 637938 584960 638028
rect 582649 637936 584960 637938
rect 582649 637880 582654 637936
rect 582710 637880 584960 637936
rect 582649 637878 584960 637880
rect 582649 637875 582715 637878
rect 583520 637788 584960 637878
rect -960 637108 480 637348
rect 580165 633858 580231 633861
rect 583520 633858 584960 633948
rect 580165 633856 584960 633858
rect 580165 633800 580170 633856
rect 580226 633800 584960 633856
rect 580165 633798 584960 633800
rect 580165 633795 580231 633798
rect 583520 633708 584960 633798
rect -960 633028 480 633268
rect 580165 629778 580231 629781
rect 583520 629778 584960 629868
rect 580165 629776 584960 629778
rect 580165 629720 580170 629776
rect 580226 629720 584960 629776
rect 580165 629718 584960 629720
rect 580165 629715 580231 629718
rect 583520 629628 584960 629718
rect -960 629098 480 629188
rect 3417 629098 3483 629101
rect -960 629096 3483 629098
rect -960 629040 3422 629096
rect 3478 629040 3483 629096
rect -960 629038 3483 629040
rect -960 628948 480 629038
rect 3417 629035 3483 629038
rect 580533 625698 580599 625701
rect 583520 625698 584960 625788
rect 580533 625696 584960 625698
rect 580533 625640 580538 625696
rect 580594 625640 584960 625696
rect 580533 625638 584960 625640
rect 580533 625635 580599 625638
rect 583520 625548 584960 625638
rect -960 625018 480 625108
rect 3233 625018 3299 625021
rect -960 625016 3299 625018
rect -960 624960 3238 625016
rect 3294 624960 3299 625016
rect -960 624958 3299 624960
rect -960 624868 480 624958
rect 3233 624955 3299 624958
rect 582557 621618 582623 621621
rect 583520 621618 584960 621708
rect 582557 621616 584960 621618
rect 582557 621560 582562 621616
rect 582618 621560 584960 621616
rect 582557 621558 584960 621560
rect 582557 621555 582623 621558
rect 583520 621468 584960 621558
rect -960 620938 480 621028
rect 3417 620938 3483 620941
rect -960 620936 3483 620938
rect -960 620880 3422 620936
rect 3478 620880 3483 620936
rect -960 620878 3483 620880
rect -960 620788 480 620878
rect 3417 620875 3483 620878
rect 582833 617538 582899 617541
rect 583520 617538 584960 617628
rect 582833 617536 584960 617538
rect 582833 617480 582838 617536
rect 582894 617480 584960 617536
rect 582833 617478 584960 617480
rect 582833 617475 582899 617478
rect 583520 617388 584960 617478
rect -960 616858 480 616948
rect 3233 616858 3299 616861
rect -960 616856 3299 616858
rect -960 616800 3238 616856
rect 3294 616800 3299 616856
rect -960 616798 3299 616800
rect -960 616708 480 616798
rect 3233 616795 3299 616798
rect 582741 613458 582807 613461
rect 583520 613458 584960 613548
rect 582741 613456 584960 613458
rect 582741 613400 582746 613456
rect 582802 613400 584960 613456
rect 582741 613398 584960 613400
rect 582741 613395 582807 613398
rect 583520 613308 584960 613398
rect -960 612778 480 612868
rect 3417 612778 3483 612781
rect -960 612776 3483 612778
rect -960 612720 3422 612776
rect 3478 612720 3483 612776
rect -960 612718 3483 612720
rect -960 612628 480 612718
rect 3417 612715 3483 612718
rect 580165 609378 580231 609381
rect 583520 609378 584960 609468
rect 580165 609376 584960 609378
rect 580165 609320 580170 609376
rect 580226 609320 584960 609376
rect 580165 609318 584960 609320
rect 580165 609315 580231 609318
rect 583520 609228 584960 609318
rect -960 608698 480 608788
rect 3417 608698 3483 608701
rect -960 608696 3483 608698
rect -960 608640 3422 608696
rect 3478 608640 3483 608696
rect -960 608638 3483 608640
rect -960 608548 480 608638
rect 3417 608635 3483 608638
rect 580349 605298 580415 605301
rect 583520 605298 584960 605388
rect 580349 605296 584960 605298
rect 580349 605240 580354 605296
rect 580410 605240 584960 605296
rect 580349 605238 584960 605240
rect 580349 605235 580415 605238
rect 583520 605148 584960 605238
rect -960 604618 480 604708
rect 3417 604618 3483 604621
rect -960 604616 3483 604618
rect -960 604560 3422 604616
rect 3478 604560 3483 604616
rect -960 604558 3483 604560
rect -960 604468 480 604558
rect 3417 604555 3483 604558
rect 583520 601068 584960 601308
rect -960 600538 480 600628
rect 3417 600538 3483 600541
rect -960 600536 3483 600538
rect -960 600480 3422 600536
rect 3478 600480 3483 600536
rect -960 600478 3483 600480
rect -960 600388 480 600478
rect 3417 600475 3483 600478
rect -960 597138 480 597228
rect 3417 597138 3483 597141
rect -960 597136 3483 597138
rect -960 597080 3422 597136
rect 3478 597080 3483 597136
rect -960 597078 3483 597080
rect -960 596988 480 597078
rect 3417 597075 3483 597078
rect 580165 597138 580231 597141
rect 583520 597138 584960 597228
rect 580165 597136 584960 597138
rect 580165 597080 580170 597136
rect 580226 597080 584960 597136
rect 580165 597078 584960 597080
rect 580165 597075 580231 597078
rect 583520 596988 584960 597078
rect -960 592908 480 593148
rect 580165 593058 580231 593061
rect 583520 593058 584960 593148
rect 580165 593056 584960 593058
rect 580165 593000 580170 593056
rect 580226 593000 584960 593056
rect 580165 592998 584960 593000
rect 580165 592995 580231 592998
rect 583520 592908 584960 592998
rect -960 588978 480 589068
rect 3417 588978 3483 588981
rect -960 588976 3483 588978
rect -960 588920 3422 588976
rect 3478 588920 3483 588976
rect -960 588918 3483 588920
rect -960 588828 480 588918
rect 3417 588915 3483 588918
rect 580533 588978 580599 588981
rect 583520 588978 584960 589068
rect 580533 588976 584960 588978
rect 580533 588920 580538 588976
rect 580594 588920 584960 588976
rect 580533 588918 584960 588920
rect 580533 588915 580599 588918
rect 583520 588828 584960 588918
rect -960 584898 480 584988
rect 3417 584898 3483 584901
rect -960 584896 3483 584898
rect -960 584840 3422 584896
rect 3478 584840 3483 584896
rect -960 584838 3483 584840
rect -960 584748 480 584838
rect 3417 584835 3483 584838
rect 580165 584898 580231 584901
rect 583520 584898 584960 584988
rect 580165 584896 584960 584898
rect 580165 584840 580170 584896
rect 580226 584840 584960 584896
rect 580165 584838 584960 584840
rect 580165 584835 580231 584838
rect 583520 584748 584960 584838
rect 583520 581348 584960 581588
rect -960 580818 480 580908
rect 3417 580818 3483 580821
rect -960 580816 3483 580818
rect -960 580760 3422 580816
rect 3478 580760 3483 580816
rect -960 580758 3483 580760
rect -960 580668 480 580758
rect 3417 580755 3483 580758
rect 578877 577418 578943 577421
rect 583520 577418 584960 577508
rect 578877 577416 584960 577418
rect 578877 577360 578882 577416
rect 578938 577360 584960 577416
rect 578877 577358 584960 577360
rect 578877 577355 578943 577358
rect 583520 577268 584960 577358
rect -960 576738 480 576828
rect 3233 576738 3299 576741
rect -960 576736 3299 576738
rect -960 576680 3238 576736
rect 3294 576680 3299 576736
rect -960 576678 3299 576680
rect -960 576588 480 576678
rect 3233 576675 3299 576678
rect 580165 573338 580231 573341
rect 583520 573338 584960 573428
rect 580165 573336 584960 573338
rect 580165 573280 580170 573336
rect 580226 573280 584960 573336
rect 580165 573278 584960 573280
rect 580165 573275 580231 573278
rect 583520 573188 584960 573278
rect -960 572658 480 572748
rect 3417 572658 3483 572661
rect -960 572656 3483 572658
rect -960 572600 3422 572656
rect 3478 572600 3483 572656
rect -960 572598 3483 572600
rect -960 572508 480 572598
rect 3417 572595 3483 572598
rect 579705 569258 579771 569261
rect 583520 569258 584960 569348
rect 579705 569256 584960 569258
rect 579705 569200 579710 569256
rect 579766 569200 584960 569256
rect 579705 569198 584960 569200
rect 579705 569195 579771 569198
rect 583520 569108 584960 569198
rect -960 568578 480 568668
rect 3233 568578 3299 568581
rect -960 568576 3299 568578
rect -960 568520 3238 568576
rect 3294 568520 3299 568576
rect -960 568518 3299 568520
rect -960 568428 480 568518
rect 3233 568515 3299 568518
rect 580165 565178 580231 565181
rect 583520 565178 584960 565268
rect 580165 565176 584960 565178
rect 580165 565120 580170 565176
rect 580226 565120 584960 565176
rect 580165 565118 584960 565120
rect 580165 565115 580231 565118
rect 583520 565028 584960 565118
rect -960 564498 480 564588
rect 3417 564498 3483 564501
rect -960 564496 3483 564498
rect -960 564440 3422 564496
rect 3478 564440 3483 564496
rect -960 564438 3483 564440
rect -960 564348 480 564438
rect 3417 564435 3483 564438
rect 579613 561098 579679 561101
rect 583520 561098 584960 561188
rect 579613 561096 584960 561098
rect 579613 561040 579618 561096
rect 579674 561040 584960 561096
rect 579613 561038 584960 561040
rect 579613 561035 579679 561038
rect 583520 560948 584960 561038
rect -960 560418 480 560508
rect 3417 560418 3483 560421
rect -960 560416 3483 560418
rect -960 560360 3422 560416
rect 3478 560360 3483 560416
rect -960 560358 3483 560360
rect -960 560268 480 560358
rect 3417 560355 3483 560358
rect 582925 557018 582991 557021
rect 583520 557018 584960 557108
rect 582925 557016 584960 557018
rect 582925 556960 582930 557016
rect 582986 556960 584960 557016
rect 582925 556958 584960 556960
rect 582925 556955 582991 556958
rect 583520 556868 584960 556958
rect -960 556338 480 556428
rect 3417 556338 3483 556341
rect -960 556336 3483 556338
rect -960 556280 3422 556336
rect 3478 556280 3483 556336
rect -960 556278 3483 556280
rect -960 556188 480 556278
rect 3417 556275 3483 556278
rect 583520 552788 584960 553028
rect -960 552258 480 552348
rect 3417 552258 3483 552261
rect -960 552256 3483 552258
rect -960 552200 3422 552256
rect 3478 552200 3483 552256
rect -960 552198 3483 552200
rect -960 552108 480 552198
rect 3417 552195 3483 552198
rect 580073 548858 580139 548861
rect 583520 548858 584960 548948
rect 580073 548856 584960 548858
rect 580073 548800 580078 548856
rect 580134 548800 584960 548856
rect 580073 548798 584960 548800
rect 580073 548795 580139 548798
rect 583520 548708 584960 548798
rect -960 548178 480 548268
rect 3233 548178 3299 548181
rect -960 548176 3299 548178
rect -960 548120 3238 548176
rect 3294 548120 3299 548176
rect -960 548118 3299 548120
rect -960 548028 480 548118
rect 3233 548115 3299 548118
rect 580165 544778 580231 544781
rect 583520 544778 584960 544868
rect 580165 544776 584960 544778
rect 580165 544720 580170 544776
rect 580226 544720 584960 544776
rect 580165 544718 584960 544720
rect 580165 544715 580231 544718
rect 583520 544628 584960 544718
rect -960 544098 480 544188
rect 3325 544098 3391 544101
rect -960 544096 3391 544098
rect -960 544040 3330 544096
rect 3386 544040 3391 544096
rect -960 544038 3391 544040
rect -960 543948 480 544038
rect 3325 544035 3391 544038
rect 579705 540698 579771 540701
rect 583520 540698 584960 540788
rect 579705 540696 584960 540698
rect 579705 540640 579710 540696
rect 579766 540640 584960 540696
rect 579705 540638 584960 540640
rect 579705 540635 579771 540638
rect 583520 540548 584960 540638
rect -960 540018 480 540108
rect 3417 540018 3483 540021
rect -960 540016 3483 540018
rect -960 539960 3422 540016
rect 3478 539960 3483 540016
rect -960 539958 3483 539960
rect -960 539868 480 539958
rect 3417 539955 3483 539958
rect -960 536468 480 536708
rect 580165 536618 580231 536621
rect 583520 536618 584960 536708
rect 580165 536616 584960 536618
rect 580165 536560 580170 536616
rect 580226 536560 584960 536616
rect 580165 536558 584960 536560
rect 580165 536555 580231 536558
rect 583520 536468 584960 536558
rect -960 532538 480 532628
rect 3233 532538 3299 532541
rect -960 532536 3299 532538
rect -960 532480 3238 532536
rect 3294 532480 3299 532536
rect -960 532478 3299 532480
rect -960 532388 480 532478
rect 3233 532475 3299 532478
rect 583017 532538 583083 532541
rect 583520 532538 584960 532628
rect 583017 532536 584960 532538
rect 583017 532480 583022 532536
rect 583078 532480 584960 532536
rect 583017 532478 584960 532480
rect 583017 532475 583083 532478
rect 583520 532388 584960 532478
rect -960 528458 480 528548
rect 3417 528458 3483 528461
rect -960 528456 3483 528458
rect -960 528400 3422 528456
rect 3478 528400 3483 528456
rect -960 528398 3483 528400
rect -960 528308 480 528398
rect 3417 528395 3483 528398
rect 580165 528458 580231 528461
rect 583520 528458 584960 528548
rect 580165 528456 584960 528458
rect 580165 528400 580170 528456
rect 580226 528400 584960 528456
rect 580165 528398 584960 528400
rect 580165 528395 580231 528398
rect 583520 528308 584960 528398
rect -960 524378 480 524468
rect 3233 524378 3299 524381
rect -960 524376 3299 524378
rect -960 524320 3238 524376
rect 3294 524320 3299 524376
rect -960 524318 3299 524320
rect -960 524228 480 524318
rect 3233 524315 3299 524318
rect 580165 524378 580231 524381
rect 583520 524378 584960 524468
rect 580165 524376 584960 524378
rect 580165 524320 580170 524376
rect 580226 524320 584960 524376
rect 580165 524318 584960 524320
rect 580165 524315 580231 524318
rect 583520 524228 584960 524318
rect 579705 520978 579771 520981
rect 583520 520978 584960 521068
rect 579705 520976 584960 520978
rect 579705 520920 579710 520976
rect 579766 520920 584960 520976
rect 579705 520918 584960 520920
rect 579705 520915 579771 520918
rect 583520 520828 584960 520918
rect -960 520298 480 520388
rect 3417 520298 3483 520301
rect -960 520296 3483 520298
rect -960 520240 3422 520296
rect 3478 520240 3483 520296
rect -960 520238 3483 520240
rect -960 520148 480 520238
rect 3417 520235 3483 520238
rect 580165 516898 580231 516901
rect 583520 516898 584960 516988
rect 580165 516896 584960 516898
rect 580165 516840 580170 516896
rect 580226 516840 584960 516896
rect 580165 516838 584960 516840
rect 580165 516835 580231 516838
rect 583520 516748 584960 516838
rect -960 516218 480 516308
rect 3417 516218 3483 516221
rect -960 516216 3483 516218
rect -960 516160 3422 516216
rect 3478 516160 3483 516216
rect -960 516158 3483 516160
rect -960 516068 480 516158
rect 3417 516155 3483 516158
rect 579613 512818 579679 512821
rect 583520 512818 584960 512908
rect 579613 512816 584960 512818
rect 579613 512760 579618 512816
rect 579674 512760 584960 512816
rect 579613 512758 584960 512760
rect 579613 512755 579679 512758
rect 583520 512668 584960 512758
rect -960 512138 480 512228
rect 3417 512138 3483 512141
rect -960 512136 3483 512138
rect -960 512080 3422 512136
rect 3478 512080 3483 512136
rect -960 512078 3483 512080
rect -960 511988 480 512078
rect 3417 512075 3483 512078
rect 580165 508738 580231 508741
rect 583520 508738 584960 508828
rect 580165 508736 584960 508738
rect 580165 508680 580170 508736
rect 580226 508680 584960 508736
rect 580165 508678 584960 508680
rect 580165 508675 580231 508678
rect 583520 508588 584960 508678
rect -960 508058 480 508148
rect 3417 508058 3483 508061
rect -960 508056 3483 508058
rect -960 508000 3422 508056
rect 3478 508000 3483 508056
rect -960 507998 3483 508000
rect -960 507908 480 507998
rect 3417 507995 3483 507998
rect 580073 504658 580139 504661
rect 583520 504658 584960 504748
rect 580073 504656 584960 504658
rect 580073 504600 580078 504656
rect 580134 504600 584960 504656
rect 580073 504598 584960 504600
rect 580073 504595 580139 504598
rect 583520 504508 584960 504598
rect -960 503978 480 504068
rect 3233 503978 3299 503981
rect -960 503976 3299 503978
rect -960 503920 3238 503976
rect 3294 503920 3299 503976
rect -960 503918 3299 503920
rect -960 503828 480 503918
rect 3233 503915 3299 503918
rect 580165 500578 580231 500581
rect 583520 500578 584960 500668
rect 580165 500576 584960 500578
rect 580165 500520 580170 500576
rect 580226 500520 584960 500576
rect 580165 500518 584960 500520
rect 580165 500515 580231 500518
rect 583520 500428 584960 500518
rect -960 499898 480 499988
rect 3325 499898 3391 499901
rect -960 499896 3391 499898
rect -960 499840 3330 499896
rect 3386 499840 3391 499896
rect -960 499838 3391 499840
rect -960 499748 480 499838
rect 3325 499835 3391 499838
rect 580165 496498 580231 496501
rect 583520 496498 584960 496588
rect 580165 496496 584960 496498
rect 580165 496440 580170 496496
rect 580226 496440 584960 496496
rect 580165 496438 584960 496440
rect 580165 496435 580231 496438
rect 583520 496348 584960 496438
rect -960 495818 480 495908
rect 2865 495818 2931 495821
rect -960 495816 2931 495818
rect -960 495760 2870 495816
rect 2926 495760 2931 495816
rect -960 495758 2931 495760
rect -960 495668 480 495758
rect 2865 495755 2931 495758
rect 583520 492268 584960 492508
rect -960 491738 480 491828
rect 3417 491738 3483 491741
rect -960 491736 3483 491738
rect -960 491680 3422 491736
rect 3478 491680 3483 491736
rect -960 491678 3483 491680
rect -960 491588 480 491678
rect 3417 491675 3483 491678
rect 580165 488338 580231 488341
rect 583520 488338 584960 488428
rect 580165 488336 584960 488338
rect 580165 488280 580170 488336
rect 580226 488280 584960 488336
rect 580165 488278 584960 488280
rect 580165 488275 580231 488278
rect 583520 488188 584960 488278
rect -960 487658 480 487748
rect 3417 487658 3483 487661
rect -960 487656 3483 487658
rect -960 487600 3422 487656
rect 3478 487600 3483 487656
rect -960 487598 3483 487600
rect -960 487508 480 487598
rect 3417 487595 3483 487598
rect 580165 484258 580231 484261
rect 583520 484258 584960 484348
rect 580165 484256 584960 484258
rect 580165 484200 580170 484256
rect 580226 484200 584960 484256
rect 580165 484198 584960 484200
rect 580165 484195 580231 484198
rect 583520 484108 584960 484198
rect -960 483578 480 483668
rect 3509 483578 3575 483581
rect -960 483576 3575 483578
rect -960 483520 3514 483576
rect 3570 483520 3575 483576
rect -960 483518 3575 483520
rect -960 483428 480 483518
rect 3509 483515 3575 483518
rect -960 480178 480 480268
rect 3417 480178 3483 480181
rect -960 480176 3483 480178
rect -960 480120 3422 480176
rect 3478 480120 3483 480176
rect -960 480118 3483 480120
rect -960 480028 480 480118
rect 3417 480115 3483 480118
rect 580165 480178 580231 480181
rect 583520 480178 584960 480268
rect 580165 480176 584960 480178
rect 580165 480120 580170 480176
rect 580226 480120 584960 480176
rect 580165 480118 584960 480120
rect 580165 480115 580231 480118
rect 583520 480028 584960 480118
rect -960 476098 480 476188
rect 3233 476098 3299 476101
rect -960 476096 3299 476098
rect -960 476040 3238 476096
rect 3294 476040 3299 476096
rect -960 476038 3299 476040
rect -960 475948 480 476038
rect 3233 476035 3299 476038
rect 580165 476098 580231 476101
rect 583520 476098 584960 476188
rect 580165 476096 584960 476098
rect 580165 476040 580170 476096
rect 580226 476040 584960 476096
rect 580165 476038 584960 476040
rect 580165 476035 580231 476038
rect 583520 475948 584960 476038
rect -960 472018 480 472108
rect 3417 472018 3483 472021
rect -960 472016 3483 472018
rect -960 471960 3422 472016
rect 3478 471960 3483 472016
rect -960 471958 3483 471960
rect -960 471868 480 471958
rect 3417 471955 3483 471958
rect 580165 472018 580231 472021
rect 583520 472018 584960 472108
rect 580165 472016 584960 472018
rect 580165 471960 580170 472016
rect 580226 471960 584960 472016
rect 580165 471958 584960 471960
rect 580165 471955 580231 471958
rect 583520 471868 584960 471958
rect -960 467938 480 468028
rect 3417 467938 3483 467941
rect -960 467936 3483 467938
rect -960 467880 3422 467936
rect 3478 467880 3483 467936
rect -960 467878 3483 467880
rect -960 467788 480 467878
rect 3417 467875 3483 467878
rect 580165 467938 580231 467941
rect 583520 467938 584960 468028
rect 580165 467936 584960 467938
rect 580165 467880 580170 467936
rect 580226 467880 584960 467936
rect 580165 467878 584960 467880
rect 580165 467875 580231 467878
rect 583520 467788 584960 467878
rect -960 463858 480 463948
rect 3417 463858 3483 463861
rect -960 463856 3483 463858
rect -960 463800 3422 463856
rect 3478 463800 3483 463856
rect -960 463798 3483 463800
rect -960 463708 480 463798
rect 3417 463795 3483 463798
rect 580165 463858 580231 463861
rect 583520 463858 584960 463948
rect 580165 463856 584960 463858
rect 580165 463800 580170 463856
rect 580226 463800 584960 463856
rect 580165 463798 584960 463800
rect 580165 463795 580231 463798
rect 583520 463708 584960 463798
rect 580165 460458 580231 460461
rect 583520 460458 584960 460548
rect 580165 460456 584960 460458
rect 580165 460400 580170 460456
rect 580226 460400 584960 460456
rect 580165 460398 584960 460400
rect 580165 460395 580231 460398
rect 583520 460308 584960 460398
rect -960 459778 480 459868
rect 3417 459778 3483 459781
rect -960 459776 3483 459778
rect -960 459720 3422 459776
rect 3478 459720 3483 459776
rect -960 459718 3483 459720
rect -960 459628 480 459718
rect 3417 459715 3483 459718
rect 580073 456378 580139 456381
rect 583520 456378 584960 456468
rect 580073 456376 584960 456378
rect 580073 456320 580078 456376
rect 580134 456320 584960 456376
rect 580073 456318 584960 456320
rect 580073 456315 580139 456318
rect 583520 456228 584960 456318
rect -960 455698 480 455788
rect 3233 455698 3299 455701
rect -960 455696 3299 455698
rect -960 455640 3238 455696
rect 3294 455640 3299 455696
rect -960 455638 3299 455640
rect -960 455548 480 455638
rect 3233 455635 3299 455638
rect 580165 452298 580231 452301
rect 583520 452298 584960 452388
rect 580165 452296 584960 452298
rect 580165 452240 580170 452296
rect 580226 452240 584960 452296
rect 580165 452238 584960 452240
rect 580165 452235 580231 452238
rect 583520 452148 584960 452238
rect -960 451618 480 451708
rect 3325 451618 3391 451621
rect -960 451616 3391 451618
rect -960 451560 3330 451616
rect 3386 451560 3391 451616
rect -960 451558 3391 451560
rect -960 451468 480 451558
rect 3325 451555 3391 451558
rect 579705 448218 579771 448221
rect 583520 448218 584960 448308
rect 579705 448216 584960 448218
rect 579705 448160 579710 448216
rect 579766 448160 584960 448216
rect 579705 448158 584960 448160
rect 579705 448155 579771 448158
rect 583520 448068 584960 448158
rect -960 447388 480 447628
rect 580165 444138 580231 444141
rect 583520 444138 584960 444228
rect 580165 444136 584960 444138
rect 580165 444080 580170 444136
rect 580226 444080 584960 444136
rect 580165 444078 584960 444080
rect 580165 444075 580231 444078
rect 583520 443988 584960 444078
rect -960 443458 480 443548
rect 3417 443458 3483 443461
rect -960 443456 3483 443458
rect -960 443400 3422 443456
rect 3478 443400 3483 443456
rect -960 443398 3483 443400
rect -960 443308 480 443398
rect 3417 443395 3483 443398
rect 581821 440058 581887 440061
rect 583520 440058 584960 440148
rect 581821 440056 584960 440058
rect 581821 440000 581826 440056
rect 581882 440000 584960 440056
rect 581821 439998 584960 440000
rect 581821 439995 581887 439998
rect 583520 439908 584960 439998
rect -960 439378 480 439468
rect 3417 439378 3483 439381
rect -960 439376 3483 439378
rect -960 439320 3422 439376
rect 3478 439320 3483 439376
rect -960 439318 3483 439320
rect -960 439228 480 439318
rect 3417 439315 3483 439318
rect 580165 435978 580231 435981
rect 583520 435978 584960 436068
rect 580165 435976 584960 435978
rect 580165 435920 580170 435976
rect 580226 435920 584960 435976
rect 580165 435918 584960 435920
rect 580165 435915 580231 435918
rect 583520 435828 584960 435918
rect -960 435148 480 435388
rect 580165 431898 580231 431901
rect 583520 431898 584960 431988
rect 580165 431896 584960 431898
rect 580165 431840 580170 431896
rect 580226 431840 584960 431896
rect 580165 431838 584960 431840
rect 580165 431835 580231 431838
rect 583520 431748 584960 431838
rect -960 431218 480 431308
rect 3509 431218 3575 431221
rect -960 431216 3575 431218
rect -960 431160 3514 431216
rect 3570 431160 3575 431216
rect -960 431158 3575 431160
rect -960 431068 480 431158
rect 3509 431155 3575 431158
rect 580165 427818 580231 427821
rect 583520 427818 584960 427908
rect 580165 427816 584960 427818
rect 580165 427760 580170 427816
rect 580226 427760 584960 427816
rect 580165 427758 584960 427760
rect 580165 427755 580231 427758
rect 583520 427668 584960 427758
rect -960 427138 480 427228
rect 2865 427138 2931 427141
rect -960 427136 2931 427138
rect -960 427080 2870 427136
rect 2926 427080 2931 427136
rect -960 427078 2931 427080
rect -960 426988 480 427078
rect 2865 427075 2931 427078
rect 580165 423738 580231 423741
rect 583520 423738 584960 423828
rect 580165 423736 584960 423738
rect 580165 423680 580170 423736
rect 580226 423680 584960 423736
rect 580165 423678 584960 423680
rect 580165 423675 580231 423678
rect 583520 423588 584960 423678
rect -960 423058 480 423148
rect 2957 423058 3023 423061
rect -960 423056 3023 423058
rect -960 423000 2962 423056
rect 3018 423000 3023 423056
rect -960 422998 3023 423000
rect -960 422908 480 422998
rect 2957 422995 3023 422998
rect -960 419658 480 419748
rect 3509 419658 3575 419661
rect -960 419656 3575 419658
rect -960 419600 3514 419656
rect 3570 419600 3575 419656
rect -960 419598 3575 419600
rect -960 419508 480 419598
rect 3509 419595 3575 419598
rect 580165 419658 580231 419661
rect 583520 419658 584960 419748
rect 580165 419656 584960 419658
rect 580165 419600 580170 419656
rect 580226 419600 584960 419656
rect 580165 419598 584960 419600
rect 580165 419595 580231 419598
rect 583520 419508 584960 419598
rect -960 415578 480 415668
rect 3509 415578 3575 415581
rect -960 415576 3575 415578
rect -960 415520 3514 415576
rect 3570 415520 3575 415576
rect -960 415518 3575 415520
rect -960 415428 480 415518
rect 3509 415515 3575 415518
rect 580165 415578 580231 415581
rect 583520 415578 584960 415668
rect 580165 415576 584960 415578
rect 580165 415520 580170 415576
rect 580226 415520 584960 415576
rect 580165 415518 584960 415520
rect 580165 415515 580231 415518
rect 583520 415428 584960 415518
rect -960 411498 480 411588
rect 3509 411498 3575 411501
rect -960 411496 3575 411498
rect -960 411440 3514 411496
rect 3570 411440 3575 411496
rect -960 411438 3575 411440
rect -960 411348 480 411438
rect 3509 411435 3575 411438
rect 579981 411498 580047 411501
rect 583520 411498 584960 411588
rect 579981 411496 584960 411498
rect 579981 411440 579986 411496
rect 580042 411440 584960 411496
rect 579981 411438 584960 411440
rect 579981 411435 580047 411438
rect 583520 411348 584960 411438
rect -960 407418 480 407508
rect 3509 407418 3575 407421
rect -960 407416 3575 407418
rect -960 407360 3514 407416
rect 3570 407360 3575 407416
rect -960 407358 3575 407360
rect -960 407268 480 407358
rect 3509 407355 3575 407358
rect 580165 407418 580231 407421
rect 583520 407418 584960 407508
rect 580165 407416 584960 407418
rect 580165 407360 580170 407416
rect 580226 407360 584960 407416
rect 580165 407358 584960 407360
rect 580165 407355 580231 407358
rect 583520 407268 584960 407358
rect 580165 404018 580231 404021
rect 583520 404018 584960 404108
rect 580165 404016 584960 404018
rect 580165 403960 580170 404016
rect 580226 403960 584960 404016
rect 580165 403958 584960 403960
rect 580165 403955 580231 403958
rect 583520 403868 584960 403958
rect -960 403338 480 403428
rect 3325 403338 3391 403341
rect -960 403336 3391 403338
rect -960 403280 3330 403336
rect 3386 403280 3391 403336
rect -960 403278 3391 403280
rect -960 403188 480 403278
rect 3325 403275 3391 403278
rect 579705 399938 579771 399941
rect 583520 399938 584960 400028
rect 579705 399936 584960 399938
rect 579705 399880 579710 399936
rect 579766 399880 584960 399936
rect 579705 399878 584960 399880
rect 579705 399875 579771 399878
rect 583520 399788 584960 399878
rect -960 399108 480 399348
rect 580165 395858 580231 395861
rect 583520 395858 584960 395948
rect 580165 395856 584960 395858
rect 580165 395800 580170 395856
rect 580226 395800 584960 395856
rect 580165 395798 584960 395800
rect 580165 395795 580231 395798
rect 583520 395708 584960 395798
rect -960 395028 480 395268
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect -960 391098 480 391188
rect 3509 391098 3575 391101
rect -960 391096 3575 391098
rect -960 391040 3514 391096
rect 3570 391040 3575 391096
rect -960 391038 3575 391040
rect -960 390948 480 391038
rect 3509 391035 3575 391038
rect 580165 387698 580231 387701
rect 583520 387698 584960 387788
rect 580165 387696 584960 387698
rect 580165 387640 580170 387696
rect 580226 387640 584960 387696
rect 580165 387638 584960 387640
rect 580165 387635 580231 387638
rect 583520 387548 584960 387638
rect -960 387018 480 387108
rect 3509 387018 3575 387021
rect -960 387016 3575 387018
rect -960 386960 3514 387016
rect 3570 386960 3575 387016
rect -960 386958 3575 386960
rect -960 386868 480 386958
rect 3509 386955 3575 386958
rect 578969 383618 579035 383621
rect 583520 383618 584960 383708
rect 578969 383616 584960 383618
rect 578969 383560 578974 383616
rect 579030 383560 584960 383616
rect 578969 383558 584960 383560
rect 578969 383555 579035 383558
rect 583520 383468 584960 383558
rect -960 382788 480 383028
rect 580441 379538 580507 379541
rect 583520 379538 584960 379628
rect 580441 379536 584960 379538
rect 580441 379480 580446 379536
rect 580502 379480 584960 379536
rect 580441 379478 584960 379480
rect 580441 379475 580507 379478
rect 583520 379388 584960 379478
rect -960 378858 480 378948
rect 2865 378858 2931 378861
rect -960 378856 2931 378858
rect -960 378800 2870 378856
rect 2926 378800 2931 378856
rect -960 378798 2931 378800
rect -960 378708 480 378798
rect 2865 378795 2931 378798
rect 580165 375458 580231 375461
rect 583520 375458 584960 375548
rect 580165 375456 584960 375458
rect 580165 375400 580170 375456
rect 580226 375400 584960 375456
rect 580165 375398 584960 375400
rect 580165 375395 580231 375398
rect 583520 375308 584960 375398
rect -960 374778 480 374868
rect 2957 374778 3023 374781
rect -960 374776 3023 374778
rect -960 374720 2962 374776
rect 3018 374720 3023 374776
rect -960 374718 3023 374720
rect -960 374628 480 374718
rect 2957 374715 3023 374718
rect 579797 371378 579863 371381
rect 583520 371378 584960 371468
rect 579797 371376 584960 371378
rect 579797 371320 579802 371376
rect 579858 371320 584960 371376
rect 579797 371318 584960 371320
rect 579797 371315 579863 371318
rect 583520 371228 584960 371318
rect -960 370698 480 370788
rect 3049 370698 3115 370701
rect -960 370696 3115 370698
rect -960 370640 3054 370696
rect 3110 370640 3115 370696
rect -960 370638 3115 370640
rect -960 370548 480 370638
rect 3049 370635 3115 370638
rect 580165 367298 580231 367301
rect 583520 367298 584960 367388
rect 580165 367296 584960 367298
rect 580165 367240 580170 367296
rect 580226 367240 584960 367296
rect 580165 367238 584960 367240
rect 580165 367235 580231 367238
rect 583520 367148 584960 367238
rect -960 366468 480 366708
rect 583520 363068 584960 363308
rect -960 362538 480 362628
rect 3049 362538 3115 362541
rect -960 362536 3115 362538
rect -960 362480 3054 362536
rect 3110 362480 3115 362536
rect -960 362478 3115 362480
rect -960 362388 480 362478
rect 3049 362475 3115 362478
rect -960 359138 480 359228
rect 3325 359138 3391 359141
rect -960 359136 3391 359138
rect -960 359080 3330 359136
rect 3386 359080 3391 359136
rect -960 359078 3391 359080
rect -960 358988 480 359078
rect 3325 359075 3391 359078
rect 580165 359138 580231 359141
rect 583520 359138 584960 359228
rect 580165 359136 584960 359138
rect 580165 359080 580170 359136
rect 580226 359080 584960 359136
rect 580165 359078 584960 359080
rect 580165 359075 580231 359078
rect 583520 358988 584960 359078
rect -960 355058 480 355148
rect 3325 355058 3391 355061
rect -960 355056 3391 355058
rect -960 355000 3330 355056
rect 3386 355000 3391 355056
rect -960 354998 3391 355000
rect -960 354908 480 354998
rect 3325 354995 3391 354998
rect 580165 355058 580231 355061
rect 583520 355058 584960 355148
rect 580165 355056 584960 355058
rect 580165 355000 580170 355056
rect 580226 355000 584960 355056
rect 580165 354998 584960 355000
rect 580165 354995 580231 354998
rect 583520 354908 584960 354998
rect -960 350978 480 351068
rect 3509 350978 3575 350981
rect -960 350976 3575 350978
rect -960 350920 3514 350976
rect 3570 350920 3575 350976
rect -960 350918 3575 350920
rect -960 350828 480 350918
rect 3509 350915 3575 350918
rect 580165 350978 580231 350981
rect 583520 350978 584960 351068
rect 580165 350976 584960 350978
rect 580165 350920 580170 350976
rect 580226 350920 584960 350976
rect 580165 350918 584960 350920
rect 580165 350915 580231 350918
rect 583520 350828 584960 350918
rect -960 346898 480 346988
rect 3325 346898 3391 346901
rect -960 346896 3391 346898
rect -960 346840 3330 346896
rect 3386 346840 3391 346896
rect -960 346838 3391 346840
rect -960 346748 480 346838
rect 3325 346835 3391 346838
rect 580165 346898 580231 346901
rect 583520 346898 584960 346988
rect 580165 346896 584960 346898
rect 580165 346840 580170 346896
rect 580226 346840 584960 346896
rect 580165 346838 584960 346840
rect 580165 346835 580231 346838
rect 583520 346748 584960 346838
rect 579705 343498 579771 343501
rect 583520 343498 584960 343588
rect 579705 343496 584960 343498
rect 579705 343440 579710 343496
rect 579766 343440 584960 343496
rect 579705 343438 584960 343440
rect 579705 343435 579771 343438
rect 583520 343348 584960 343438
rect -960 342818 480 342908
rect 3509 342818 3575 342821
rect -960 342816 3575 342818
rect -960 342760 3514 342816
rect 3570 342760 3575 342816
rect -960 342758 3575 342760
rect -960 342668 480 342758
rect 3509 342755 3575 342758
rect 579613 339418 579679 339421
rect 583520 339418 584960 339508
rect 579613 339416 584960 339418
rect 579613 339360 579618 339416
rect 579674 339360 584960 339416
rect 579613 339358 584960 339360
rect 579613 339355 579679 339358
rect 583520 339268 584960 339358
rect -960 338738 480 338828
rect 3509 338738 3575 338741
rect -960 338736 3575 338738
rect -960 338680 3514 338736
rect 3570 338680 3575 338736
rect -960 338678 3575 338680
rect -960 338588 480 338678
rect 3509 338675 3575 338678
rect 583520 335188 584960 335428
rect -960 334508 480 334748
rect 579705 331258 579771 331261
rect 583520 331258 584960 331348
rect 579705 331256 584960 331258
rect 579705 331200 579710 331256
rect 579766 331200 584960 331256
rect 579705 331198 584960 331200
rect 579705 331195 579771 331198
rect 583520 331108 584960 331198
rect -960 330578 480 330668
rect 2957 330578 3023 330581
rect -960 330576 3023 330578
rect -960 330520 2962 330576
rect 3018 330520 3023 330576
rect -960 330518 3023 330520
rect -960 330428 480 330518
rect 2957 330515 3023 330518
rect 580625 327178 580691 327181
rect 583520 327178 584960 327268
rect 580625 327176 584960 327178
rect 580625 327120 580630 327176
rect 580686 327120 584960 327176
rect 580625 327118 584960 327120
rect 580625 327115 580691 327118
rect 583520 327028 584960 327118
rect -960 326348 480 326588
rect 579061 323098 579127 323101
rect 583520 323098 584960 323188
rect 579061 323096 584960 323098
rect 579061 323040 579066 323096
rect 579122 323040 584960 323096
rect 579061 323038 584960 323040
rect 579061 323035 579127 323038
rect 583520 322948 584960 323038
rect -960 322418 480 322508
rect 3049 322418 3115 322421
rect -960 322416 3115 322418
rect -960 322360 3054 322416
rect 3110 322360 3115 322416
rect -960 322358 3115 322360
rect -960 322268 480 322358
rect 3049 322355 3115 322358
rect 579705 319018 579771 319021
rect 583520 319018 584960 319108
rect 579705 319016 584960 319018
rect 579705 318960 579710 319016
rect 579766 318960 584960 319016
rect 579705 318958 584960 318960
rect 579705 318955 579771 318958
rect 583520 318868 584960 318958
rect -960 318338 480 318428
rect 3509 318338 3575 318341
rect -960 318336 3575 318338
rect -960 318280 3514 318336
rect 3570 318280 3575 318336
rect -960 318278 3575 318280
rect -960 318188 480 318278
rect 3509 318275 3575 318278
rect 579613 314938 579679 314941
rect 583520 314938 584960 315028
rect 579613 314936 584960 314938
rect 579613 314880 579618 314936
rect 579674 314880 584960 314936
rect 579613 314878 584960 314880
rect 579613 314875 579679 314878
rect 583520 314788 584960 314878
rect -960 314258 480 314348
rect 3049 314258 3115 314261
rect -960 314256 3115 314258
rect -960 314200 3054 314256
rect 3110 314200 3115 314256
rect -960 314198 3115 314200
rect -960 314108 480 314198
rect 3049 314195 3115 314198
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 310178 480 310268
rect 3141 310178 3207 310181
rect -960 310176 3207 310178
rect -960 310120 3146 310176
rect 3202 310120 3207 310176
rect -960 310118 3207 310120
rect -960 310028 480 310118
rect 3141 310115 3207 310118
rect 580165 306778 580231 306781
rect 583520 306778 584960 306868
rect 580165 306776 584960 306778
rect 580165 306720 580170 306776
rect 580226 306720 584960 306776
rect 580165 306718 584960 306720
rect 580165 306715 580231 306718
rect 583520 306628 584960 306718
rect -960 306098 480 306188
rect 3233 306098 3299 306101
rect -960 306096 3299 306098
rect -960 306040 3238 306096
rect 3294 306040 3299 306096
rect -960 306038 3299 306040
rect -960 305948 480 306038
rect 3233 306035 3299 306038
rect 580165 302698 580231 302701
rect 583520 302698 584960 302788
rect 580165 302696 584960 302698
rect 580165 302640 580170 302696
rect 580226 302640 584960 302696
rect 580165 302638 584960 302640
rect 580165 302635 580231 302638
rect 583520 302548 584960 302638
rect -960 302018 480 302108
rect 3141 302018 3207 302021
rect -960 302016 3207 302018
rect -960 301960 3146 302016
rect 3202 301960 3207 302016
rect -960 301958 3207 301960
rect -960 301868 480 301958
rect 3141 301955 3207 301958
rect -960 298618 480 298708
rect 3325 298618 3391 298621
rect -960 298616 3391 298618
rect -960 298560 3330 298616
rect 3386 298560 3391 298616
rect -960 298558 3391 298560
rect -960 298468 480 298558
rect 3325 298555 3391 298558
rect 579153 298618 579219 298621
rect 583520 298618 584960 298708
rect 579153 298616 584960 298618
rect 579153 298560 579158 298616
rect 579214 298560 584960 298616
rect 579153 298558 584960 298560
rect 579153 298555 579219 298558
rect 583520 298468 584960 298558
rect -960 294538 480 294628
rect 3509 294538 3575 294541
rect -960 294536 3575 294538
rect -960 294480 3514 294536
rect 3570 294480 3575 294536
rect -960 294478 3575 294480
rect -960 294388 480 294478
rect 3509 294475 3575 294478
rect 580165 294538 580231 294541
rect 583520 294538 584960 294628
rect 580165 294536 584960 294538
rect 580165 294480 580170 294536
rect 580226 294480 584960 294536
rect 580165 294478 584960 294480
rect 580165 294475 580231 294478
rect 583520 294388 584960 294478
rect -960 290458 480 290548
rect 3509 290458 3575 290461
rect -960 290456 3575 290458
rect -960 290400 3514 290456
rect 3570 290400 3575 290456
rect -960 290398 3575 290400
rect -960 290308 480 290398
rect 3509 290395 3575 290398
rect 579981 290458 580047 290461
rect 583520 290458 584960 290548
rect 579981 290456 584960 290458
rect 579981 290400 579986 290456
rect 580042 290400 584960 290456
rect 579981 290398 584960 290400
rect 579981 290395 580047 290398
rect 583520 290308 584960 290398
rect -960 286378 480 286468
rect 2865 286378 2931 286381
rect -960 286376 2931 286378
rect -960 286320 2870 286376
rect 2926 286320 2931 286376
rect -960 286318 2931 286320
rect -960 286228 480 286318
rect 2865 286315 2931 286318
rect 579981 286378 580047 286381
rect 583520 286378 584960 286468
rect 579981 286376 584960 286378
rect 579981 286320 579986 286376
rect 580042 286320 584960 286376
rect 579981 286318 584960 286320
rect 579981 286315 580047 286318
rect 583520 286228 584960 286318
rect 580165 282978 580231 282981
rect 583520 282978 584960 283068
rect 580165 282976 584960 282978
rect 580165 282920 580170 282976
rect 580226 282920 584960 282976
rect 580165 282918 584960 282920
rect 580165 282915 580231 282918
rect 583520 282828 584960 282918
rect -960 282298 480 282388
rect 2957 282298 3023 282301
rect -960 282296 3023 282298
rect -960 282240 2962 282296
rect 3018 282240 3023 282296
rect -960 282238 3023 282240
rect -960 282148 480 282238
rect 2957 282235 3023 282238
rect 580165 278898 580231 278901
rect 583520 278898 584960 278988
rect 580165 278896 584960 278898
rect 580165 278840 580170 278896
rect 580226 278840 584960 278896
rect 580165 278838 584960 278840
rect 580165 278835 580231 278838
rect 583520 278748 584960 278838
rect -960 278218 480 278308
rect 3049 278218 3115 278221
rect -960 278216 3115 278218
rect -960 278160 3054 278216
rect 3110 278160 3115 278216
rect -960 278158 3115 278160
rect -960 278068 480 278158
rect 3049 278155 3115 278158
rect 580165 274818 580231 274821
rect 583520 274818 584960 274908
rect 580165 274816 584960 274818
rect 580165 274760 580170 274816
rect 580226 274760 584960 274816
rect 580165 274758 584960 274760
rect 580165 274755 580231 274758
rect 583520 274668 584960 274758
rect -960 274138 480 274228
rect 3509 274138 3575 274141
rect -960 274136 3575 274138
rect -960 274080 3514 274136
rect 3570 274080 3575 274136
rect -960 274078 3575 274080
rect -960 273988 480 274078
rect 3509 274075 3575 274078
rect 579705 270738 579771 270741
rect 583520 270738 584960 270828
rect 579705 270736 584960 270738
rect 579705 270680 579710 270736
rect 579766 270680 584960 270736
rect 579705 270678 584960 270680
rect 579705 270675 579771 270678
rect 583520 270588 584960 270678
rect -960 270058 480 270148
rect 3049 270058 3115 270061
rect -960 270056 3115 270058
rect -960 270000 3054 270056
rect 3110 270000 3115 270056
rect -960 269998 3115 270000
rect -960 269908 480 269998
rect 3049 269995 3115 269998
rect 196014 269724 196020 269788
rect 196084 269786 196090 269788
rect 535453 269786 535519 269789
rect 196084 269784 535519 269786
rect 196084 269728 535458 269784
rect 535514 269728 535519 269784
rect 196084 269726 535519 269728
rect 196084 269724 196090 269726
rect 535453 269723 535519 269726
rect 194542 268364 194548 268428
rect 194612 268426 194618 268428
rect 263593 268426 263659 268429
rect 194612 268424 263659 268426
rect 194612 268368 263598 268424
rect 263654 268368 263659 268424
rect 194612 268366 263659 268368
rect 194612 268364 194618 268366
rect 263593 268363 263659 268366
rect 579613 266658 579679 266661
rect 583520 266658 584960 266748
rect 579613 266656 584960 266658
rect 579613 266600 579618 266656
rect 579674 266600 584960 266656
rect 579613 266598 584960 266600
rect 579613 266595 579679 266598
rect 583520 266508 584960 266598
rect -960 265978 480 266068
rect 3141 265978 3207 265981
rect -960 265976 3207 265978
rect -960 265920 3146 265976
rect 3202 265920 3207 265976
rect -960 265918 3207 265920
rect -960 265828 480 265918
rect 3141 265915 3207 265918
rect 38653 265570 38719 265573
rect 111742 265570 111748 265572
rect 38653 265568 111748 265570
rect 38653 265512 38658 265568
rect 38714 265512 111748 265568
rect 38653 265510 111748 265512
rect 38653 265507 38719 265510
rect 111742 265508 111748 265510
rect 111812 265508 111818 265572
rect 118550 263876 118556 263940
rect 118620 263938 118626 263940
rect 148041 263938 148107 263941
rect 118620 263936 148107 263938
rect 118620 263880 148046 263936
rect 148102 263880 148107 263936
rect 118620 263878 148107 263880
rect 118620 263876 118626 263878
rect 148041 263875 148107 263878
rect 116894 263740 116900 263804
rect 116964 263802 116970 263804
rect 135437 263802 135503 263805
rect 136541 263802 136607 263805
rect 116964 263800 136607 263802
rect 116964 263744 135442 263800
rect 135498 263744 136546 263800
rect 136602 263744 136607 263800
rect 116964 263742 136607 263744
rect 116964 263740 116970 263742
rect 135437 263739 135503 263742
rect 136541 263739 136607 263742
rect 168925 263666 168991 263669
rect 196198 263666 196204 263668
rect 168925 263664 196204 263666
rect 168925 263608 168930 263664
rect 168986 263608 196204 263664
rect 168925 263606 196204 263608
rect 168925 263603 168991 263606
rect 196198 263604 196204 263606
rect 196268 263666 196274 263668
rect 196617 263666 196683 263669
rect 196268 263664 196683 263666
rect 196268 263608 196622 263664
rect 196678 263608 196683 263664
rect 196268 263606 196683 263608
rect 196268 263604 196274 263606
rect 196617 263603 196683 263606
rect 183001 262986 183067 262989
rect 191782 262986 191788 262988
rect 183001 262984 191788 262986
rect 183001 262928 183006 262984
rect 183062 262928 191788 262984
rect 183001 262926 191788 262928
rect 183001 262923 183067 262926
rect 191782 262924 191788 262926
rect 191852 262924 191858 262988
rect 111742 262788 111748 262852
rect 111812 262850 111818 262852
rect 112846 262850 112852 262852
rect 111812 262790 112852 262850
rect 111812 262788 111818 262790
rect 112846 262788 112852 262790
rect 112916 262850 112922 262852
rect 134885 262850 134951 262853
rect 112916 262848 134951 262850
rect 112916 262792 134890 262848
rect 134946 262792 134951 262848
rect 112916 262790 134951 262792
rect 112916 262788 112922 262790
rect 134885 262787 134951 262790
rect 179413 262850 179479 262853
rect 193254 262850 193260 262852
rect 179413 262848 193260 262850
rect 179413 262792 179418 262848
rect 179474 262792 193260 262848
rect 179413 262790 193260 262792
rect 179413 262787 179479 262790
rect 193254 262788 193260 262790
rect 193324 262850 193330 262852
rect 194542 262850 194548 262852
rect 193324 262790 194548 262850
rect 193324 262788 193330 262790
rect 194542 262788 194548 262790
rect 194612 262788 194618 262852
rect 122557 262714 122623 262717
rect 520273 262714 520339 262717
rect 122557 262712 520339 262714
rect 122557 262656 122562 262712
rect 122618 262656 520278 262712
rect 520334 262656 520339 262712
rect 122557 262654 520339 262656
rect 122557 262651 122623 262654
rect 520273 262651 520339 262654
rect 185485 262578 185551 262581
rect 196014 262578 196020 262580
rect 185485 262576 196020 262578
rect 185485 262520 185490 262576
rect 185546 262520 196020 262576
rect 185485 262518 196020 262520
rect 185485 262515 185551 262518
rect 196014 262516 196020 262518
rect 196084 262516 196090 262580
rect 580257 262578 580323 262581
rect 583520 262578 584960 262668
rect 580257 262576 584960 262578
rect 580257 262520 580262 262576
rect 580318 262520 584960 262576
rect 580257 262518 584960 262520
rect 580257 262515 580323 262518
rect 181437 262442 181503 262445
rect 197486 262442 197492 262444
rect 181437 262440 197492 262442
rect 181437 262384 181442 262440
rect 181498 262384 197492 262440
rect 181437 262382 197492 262384
rect 181437 262379 181503 262382
rect 197486 262380 197492 262382
rect 197556 262380 197562 262444
rect 583520 262428 584960 262518
rect 121545 262308 121611 262309
rect 121494 262244 121500 262308
rect 121564 262306 121611 262308
rect 121564 262304 121656 262306
rect 121606 262248 121656 262304
rect 121564 262246 121656 262248
rect 121564 262244 121611 262246
rect 121545 262243 121611 262244
rect -960 261898 480 261988
rect 3049 261898 3115 261901
rect -960 261896 3115 261898
rect -960 261840 3054 261896
rect 3110 261840 3115 261896
rect -960 261838 3115 261840
rect -960 261748 480 261838
rect 3049 261835 3115 261838
rect 121310 260068 121316 260132
rect 121380 260130 121386 260132
rect 138105 260130 138171 260133
rect 121380 260128 138171 260130
rect 121380 260072 138110 260128
rect 138166 260072 138171 260128
rect 121380 260070 138171 260072
rect 121380 260068 121386 260070
rect 138105 260067 138171 260070
rect 122557 259996 122623 259997
rect 122557 259992 122604 259996
rect 122668 259994 122674 259996
rect 182173 259994 182239 259997
rect 183369 259994 183435 259997
rect 122557 259936 122562 259992
rect 122557 259932 122604 259936
rect 122668 259934 122714 259994
rect 182173 259992 183435 259994
rect 182173 259936 182178 259992
rect 182234 259936 183374 259992
rect 183430 259936 183435 259992
rect 182173 259934 183435 259936
rect 122668 259932 122674 259934
rect 122557 259931 122623 259932
rect 182173 259931 182239 259934
rect 183369 259931 183435 259934
rect 184933 259994 184999 259997
rect 185853 259994 185919 259997
rect 187182 259994 187188 259996
rect 184933 259992 187188 259994
rect 184933 259936 184938 259992
rect 184994 259936 185858 259992
rect 185914 259936 187188 259992
rect 184933 259934 187188 259936
rect 184933 259931 184999 259934
rect 185853 259931 185919 259934
rect 187182 259932 187188 259934
rect 187252 259932 187258 259996
rect 111558 259660 111564 259724
rect 111628 259722 111634 259724
rect 129365 259722 129431 259725
rect 111628 259720 129431 259722
rect 111628 259664 129370 259720
rect 129426 259664 129431 259720
rect 111628 259662 129431 259664
rect 111628 259660 111634 259662
rect 129365 259659 129431 259662
rect 111374 259524 111380 259588
rect 111444 259586 111450 259588
rect 131849 259586 131915 259589
rect 111444 259584 131915 259586
rect 111444 259528 131854 259584
rect 131910 259528 131915 259584
rect 111444 259526 131915 259528
rect 111444 259524 111450 259526
rect 131849 259523 131915 259526
rect 183369 259586 183435 259589
rect 195421 259586 195487 259589
rect 183369 259584 195487 259586
rect 183369 259528 183374 259584
rect 183430 259528 195426 259584
rect 195482 259528 195487 259584
rect 183369 259526 195487 259528
rect 183369 259523 183435 259526
rect 195421 259523 195487 259526
rect 186957 259316 187023 259317
rect 186957 259312 187004 259316
rect 187068 259314 187074 259316
rect 186957 259256 186962 259312
rect 186957 259252 187004 259256
rect 187068 259254 187114 259314
rect 187068 259252 187074 259254
rect 186957 259251 187023 259252
rect 580257 258498 580323 258501
rect 583520 258498 584960 258588
rect 580257 258496 584960 258498
rect 580257 258440 580262 258496
rect 580318 258440 584960 258496
rect 580257 258438 584960 258440
rect 580257 258435 580323 258438
rect 583520 258348 584960 258438
rect -960 257818 480 257908
rect 3233 257818 3299 257821
rect -960 257816 3299 257818
rect -960 257760 3238 257816
rect 3294 257760 3299 257816
rect -960 257758 3299 257760
rect -960 257668 480 257758
rect 3233 257755 3299 257758
rect 579797 254418 579863 254421
rect 583520 254418 584960 254508
rect 579797 254416 584960 254418
rect 579797 254360 579802 254416
rect 579858 254360 584960 254416
rect 579797 254358 584960 254360
rect 579797 254355 579863 254358
rect 583520 254268 584960 254358
rect -960 253738 480 253828
rect 3141 253738 3207 253741
rect -960 253736 3207 253738
rect -960 253680 3146 253736
rect 3202 253680 3207 253736
rect -960 253678 3207 253680
rect -960 253588 480 253678
rect 3141 253675 3207 253678
rect 579981 250338 580047 250341
rect 583520 250338 584960 250428
rect 579981 250336 584960 250338
rect 579981 250280 579986 250336
rect 580042 250280 584960 250336
rect 579981 250278 584960 250280
rect 579981 250275 580047 250278
rect 583520 250188 584960 250278
rect -960 249658 480 249748
rect 3509 249658 3575 249661
rect -960 249656 3575 249658
rect -960 249600 3514 249656
rect 3570 249600 3575 249656
rect -960 249598 3575 249600
rect -960 249508 480 249598
rect 3509 249595 3575 249598
rect 583520 246258 584960 246348
rect 583342 246198 584960 246258
rect 583342 246122 583402 246198
rect 583520 246122 584960 246198
rect 583342 246108 584960 246122
rect 583342 246062 583586 246108
rect -960 245428 480 245668
rect 188286 245652 188292 245716
rect 188356 245714 188362 245716
rect 583526 245714 583586 246062
rect 188356 245654 583586 245714
rect 188356 245652 188362 245654
rect 580165 242178 580231 242181
rect 583520 242178 584960 242268
rect 580165 242176 584960 242178
rect 580165 242120 580170 242176
rect 580226 242120 584960 242176
rect 580165 242118 584960 242120
rect 580165 242115 580231 242118
rect 583520 242028 584960 242118
rect -960 241498 480 241588
rect 3325 241498 3391 241501
rect -960 241496 3391 241498
rect -960 241440 3330 241496
rect 3386 241440 3391 241496
rect -960 241438 3391 241440
rect -960 241348 480 241438
rect 3325 241435 3391 241438
rect -960 238098 480 238188
rect 580165 238098 580231 238101
rect 583520 238098 584960 238188
rect -960 238038 674 238098
rect -960 237962 480 238038
rect 614 237962 674 238038
rect 580165 238096 584960 238098
rect 580165 238040 580170 238096
rect 580226 238040 584960 238096
rect 580165 238038 584960 238040
rect 580165 238035 580231 238038
rect -960 237948 674 237962
rect 583520 237948 584960 238038
rect 246 237902 674 237948
rect 246 237418 306 237902
rect 122046 237418 122052 237420
rect 246 237358 122052 237418
rect 122046 237356 122052 237358
rect 122116 237356 122122 237420
rect -960 233868 480 234108
rect 583520 234018 584960 234108
rect 583342 233958 584960 234018
rect 583342 233882 583402 233958
rect 583520 233882 584960 233958
rect 583342 233868 584960 233882
rect 583342 233822 583586 233868
rect 186814 233276 186820 233340
rect 186884 233338 186890 233340
rect 583526 233338 583586 233822
rect 186884 233278 583586 233338
rect 186884 233276 186890 233278
rect -960 229938 480 230028
rect 3325 229938 3391 229941
rect -960 229936 3391 229938
rect -960 229880 3330 229936
rect 3386 229880 3391 229936
rect -960 229878 3391 229880
rect -960 229788 480 229878
rect 3325 229875 3391 229878
rect 580717 229938 580783 229941
rect 583520 229938 584960 230028
rect 580717 229936 584960 229938
rect 580717 229880 580722 229936
rect 580778 229880 584960 229936
rect 580717 229878 584960 229880
rect 580717 229875 580783 229878
rect 583520 229788 584960 229878
rect -960 225858 480 225948
rect 3601 225858 3667 225861
rect -960 225856 3667 225858
rect -960 225800 3606 225856
rect 3662 225800 3667 225856
rect -960 225798 3667 225800
rect -960 225708 480 225798
rect 3601 225795 3667 225798
rect 579981 225858 580047 225861
rect 583520 225858 584960 225948
rect 579981 225856 584960 225858
rect 579981 225800 579986 225856
rect 580042 225800 584960 225856
rect 579981 225798 584960 225800
rect 579981 225795 580047 225798
rect 583520 225708 584960 225798
rect 583520 222308 584960 222548
rect -960 221778 480 221868
rect 3049 221778 3115 221781
rect -960 221776 3115 221778
rect -960 221720 3054 221776
rect 3110 221720 3115 221776
rect -960 221718 3115 221720
rect -960 221628 480 221718
rect 3049 221715 3115 221718
rect 583520 218378 584960 218468
rect 567150 218318 584960 218378
rect 120625 218106 120691 218109
rect 121494 218106 121500 218108
rect 120625 218104 121500 218106
rect 120625 218048 120630 218104
rect 120686 218048 121500 218104
rect 120625 218046 121500 218048
rect 120625 218043 120691 218046
rect 121494 218044 121500 218046
rect 121564 218044 121570 218108
rect 188470 218044 188476 218108
rect 188540 218106 188546 218108
rect 567150 218106 567210 218318
rect 583520 218228 584960 218318
rect 188540 218046 567210 218106
rect 188540 218044 188546 218046
rect -960 217698 480 217788
rect -960 217638 674 217698
rect -960 217562 480 217638
rect 614 217562 674 217638
rect -960 217548 674 217562
rect 246 217502 674 217548
rect 246 217018 306 217502
rect 246 216958 6930 217018
rect 6870 216746 6930 216958
rect 122230 216746 122236 216748
rect 6870 216686 122236 216746
rect 122230 216684 122236 216686
rect 122300 216684 122306 216748
rect 580809 214298 580875 214301
rect 583520 214298 584960 214388
rect 580809 214296 584960 214298
rect 580809 214240 580814 214296
rect 580870 214240 584960 214296
rect 580809 214238 584960 214240
rect 580809 214235 580875 214238
rect 583520 214148 584960 214238
rect -960 213618 480 213708
rect -960 213558 674 213618
rect -960 213482 480 213558
rect 614 213482 674 213558
rect -960 213468 674 213482
rect 246 213422 674 213468
rect 246 212938 306 213422
rect 246 212878 6930 212938
rect 6870 212666 6930 212878
rect 122414 212666 122420 212668
rect 6870 212606 122420 212666
rect 122414 212604 122420 212606
rect 122484 212604 122490 212668
rect 580901 210218 580967 210221
rect 583520 210218 584960 210308
rect 580901 210216 584960 210218
rect 580901 210160 580906 210216
rect 580962 210160 584960 210216
rect 580901 210158 584960 210160
rect 580901 210155 580967 210158
rect 583520 210068 584960 210158
rect -960 209538 480 209628
rect 3141 209538 3207 209541
rect -960 209536 3207 209538
rect -960 209480 3146 209536
rect 3202 209480 3207 209536
rect -960 209478 3207 209480
rect -960 209388 480 209478
rect 3141 209475 3207 209478
rect 583520 205988 584960 206228
rect -960 205308 480 205548
rect 92473 202194 92539 202197
rect 107377 202194 107443 202197
rect 92473 202192 107443 202194
rect 92473 202136 92478 202192
rect 92534 202136 107382 202192
rect 107438 202136 107443 202192
rect 92473 202134 107443 202136
rect 92473 202131 92539 202134
rect 107377 202131 107443 202134
rect 583520 202058 584960 202148
rect 583342 201998 584960 202058
rect 583342 201922 583402 201998
rect 583520 201922 584960 201998
rect 583342 201908 584960 201922
rect 583342 201862 583586 201908
rect 181478 201786 181484 201788
rect 176610 201726 181484 201786
rect 107377 201514 107443 201517
rect 138606 201514 138612 201516
rect 107377 201512 138612 201514
rect -960 201378 480 201468
rect 107377 201456 107382 201512
rect 107438 201456 138612 201512
rect 107377 201454 138612 201456
rect 107377 201451 107443 201454
rect 138606 201452 138612 201454
rect 138676 201452 138682 201516
rect 160318 201452 160324 201516
rect 160388 201514 160394 201516
rect 176610 201514 176670 201726
rect 181478 201724 181484 201726
rect 181548 201786 181554 201788
rect 466453 201786 466519 201789
rect 181548 201784 466519 201786
rect 181548 201728 466458 201784
rect 466514 201728 466519 201784
rect 181548 201726 466519 201728
rect 181548 201724 181554 201726
rect 466453 201723 466519 201726
rect 160388 201454 176670 201514
rect 160388 201452 160394 201454
rect 184974 201452 184980 201516
rect 185044 201514 185050 201516
rect 583526 201514 583586 201862
rect 185044 201454 583586 201514
rect 185044 201452 185050 201454
rect 4061 201378 4127 201381
rect -960 201376 4127 201378
rect -960 201320 4066 201376
rect 4122 201320 4127 201376
rect -960 201318 4127 201320
rect -960 201228 480 201318
rect 4061 201315 4127 201318
rect 207054 201044 207060 201108
rect 207124 201106 207130 201108
rect 374637 201106 374703 201109
rect 207124 201104 374703 201106
rect 207124 201048 374642 201104
rect 374698 201048 374703 201104
rect 207124 201046 374703 201048
rect 207124 201044 207130 201046
rect 374637 201043 374703 201046
rect 118693 200970 118759 200973
rect 154246 200970 154252 200972
rect 118693 200968 154252 200970
rect 118693 200912 118698 200968
rect 118754 200912 154252 200968
rect 118693 200910 154252 200912
rect 118693 200907 118759 200910
rect 154246 200908 154252 200910
rect 154316 200908 154322 200972
rect 180190 200908 180196 200972
rect 180260 200970 180266 200972
rect 186814 200970 186820 200972
rect 180260 200910 186820 200970
rect 180260 200908 180266 200910
rect 186814 200908 186820 200910
rect 186884 200908 186890 200972
rect 205030 200908 205036 200972
rect 205100 200970 205106 200972
rect 509233 200970 509299 200973
rect 205100 200968 509299 200970
rect 205100 200912 509238 200968
rect 509294 200912 509299 200968
rect 205100 200910 509299 200912
rect 205100 200908 205106 200910
rect 509233 200907 509299 200910
rect 122230 200772 122236 200836
rect 122300 200834 122306 200836
rect 122300 200774 125978 200834
rect 122300 200772 122306 200774
rect 78029 200698 78095 200701
rect 95049 200698 95115 200701
rect 78029 200696 95115 200698
rect 78029 200640 78034 200696
rect 78090 200640 95054 200696
rect 95110 200640 95115 200696
rect 78029 200638 95115 200640
rect 78029 200635 78095 200638
rect 95049 200635 95115 200638
rect 111793 200698 111859 200701
rect 122833 200698 122899 200701
rect 111793 200696 122899 200698
rect 111793 200640 111798 200696
rect 111854 200640 122838 200696
rect 122894 200640 122899 200696
rect 111793 200638 122899 200640
rect 125918 200698 125978 200774
rect 146518 200772 146524 200836
rect 146588 200834 146594 200836
rect 188286 200834 188292 200836
rect 146588 200774 188292 200834
rect 146588 200772 146594 200774
rect 188286 200772 188292 200774
rect 188356 200772 188362 200836
rect 210918 200772 210924 200836
rect 210988 200834 210994 200836
rect 561673 200834 561739 200837
rect 210988 200832 561739 200834
rect 210988 200776 561678 200832
rect 561734 200776 561739 200832
rect 210988 200774 561739 200776
rect 210988 200772 210994 200774
rect 561673 200771 561739 200774
rect 128997 200698 129063 200701
rect 125918 200696 129063 200698
rect 125918 200640 129002 200696
rect 129058 200640 129063 200696
rect 125918 200638 129063 200640
rect 111793 200635 111859 200638
rect 122833 200635 122899 200638
rect 128997 200635 129063 200638
rect 137870 200636 137876 200700
rect 137940 200698 137946 200700
rect 191189 200698 191255 200701
rect 137940 200696 191255 200698
rect 137940 200640 191194 200696
rect 191250 200640 191255 200696
rect 137940 200638 191255 200640
rect 137940 200636 137946 200638
rect 191189 200635 191255 200638
rect 211102 200636 211108 200700
rect 211172 200698 211178 200700
rect 582649 200698 582715 200701
rect 211172 200696 582715 200698
rect 211172 200640 582654 200696
rect 582710 200640 582715 200696
rect 211172 200638 582715 200640
rect 211172 200636 211178 200638
rect 582649 200635 582715 200638
rect 173566 200500 173572 200564
rect 173636 200562 173642 200564
rect 205030 200562 205036 200564
rect 173636 200502 205036 200562
rect 173636 200500 173642 200502
rect 205030 200500 205036 200502
rect 205100 200500 205106 200564
rect 122046 200364 122052 200428
rect 122116 200426 122122 200428
rect 123201 200426 123267 200429
rect 122116 200424 123267 200426
rect 122116 200368 123206 200424
rect 123262 200368 123267 200424
rect 122116 200366 123267 200368
rect 122116 200364 122122 200366
rect 123201 200363 123267 200366
rect 131481 200426 131547 200429
rect 131481 200424 140790 200426
rect 131481 200368 131486 200424
rect 131542 200368 140790 200424
rect 131481 200366 140790 200368
rect 131481 200363 131547 200366
rect 105629 200290 105695 200293
rect 132033 200290 132099 200293
rect 105629 200288 132099 200290
rect 105629 200232 105634 200288
rect 105690 200232 132038 200288
rect 132094 200232 132099 200288
rect 105629 200230 132099 200232
rect 105629 200227 105695 200230
rect 132033 200227 132099 200230
rect 132217 200290 132283 200293
rect 140446 200290 140452 200292
rect 132217 200288 140452 200290
rect 132217 200232 132222 200288
rect 132278 200232 140452 200288
rect 132217 200230 140452 200232
rect 132217 200227 132283 200230
rect 140446 200228 140452 200230
rect 140516 200228 140522 200292
rect 140730 200290 140790 200366
rect 170622 200364 170628 200428
rect 170692 200426 170698 200428
rect 178769 200426 178835 200429
rect 207054 200426 207060 200428
rect 170692 200366 177728 200426
rect 170692 200364 170698 200366
rect 158110 200290 158116 200292
rect 140730 200230 158116 200290
rect 158110 200228 158116 200230
rect 158180 200228 158186 200292
rect 160870 200228 160876 200292
rect 160940 200290 160946 200292
rect 169518 200290 169524 200292
rect 160940 200230 169524 200290
rect 160940 200228 160946 200230
rect 169518 200228 169524 200230
rect 169588 200228 169594 200292
rect 177668 200290 177728 200366
rect 178769 200424 207060 200426
rect 178769 200368 178774 200424
rect 178830 200368 207060 200424
rect 178769 200366 207060 200368
rect 178769 200363 178835 200366
rect 207054 200364 207060 200366
rect 207124 200364 207130 200428
rect 177941 200290 178007 200293
rect 177668 200288 178007 200290
rect 177668 200232 177946 200288
rect 178002 200232 178007 200288
rect 177668 200230 178007 200232
rect 177941 200227 178007 200230
rect 180425 200290 180491 200293
rect 211102 200290 211108 200292
rect 180425 200288 211108 200290
rect 180425 200232 180430 200288
rect 180486 200232 211108 200288
rect 180425 200230 211108 200232
rect 180425 200227 180491 200230
rect 211102 200228 211108 200230
rect 211172 200228 211178 200292
rect 95049 200154 95115 200157
rect 131481 200154 131547 200157
rect 95049 200152 131547 200154
rect 95049 200096 95054 200152
rect 95110 200096 131486 200152
rect 131542 200096 131547 200152
rect 95049 200094 131547 200096
rect 95049 200091 95115 200094
rect 131481 200091 131547 200094
rect 131665 200154 131731 200157
rect 152590 200154 152596 200156
rect 131665 200152 148932 200154
rect 131665 200096 131670 200152
rect 131726 200096 148932 200152
rect 131665 200094 148932 200096
rect 131665 200091 131731 200094
rect 131849 200018 131915 200021
rect 128310 200016 131915 200018
rect 128310 199960 131854 200016
rect 131910 199960 131915 200016
rect 128310 199958 131915 199960
rect 127157 199882 127223 199885
rect 128310 199882 128370 199958
rect 131849 199955 131915 199958
rect 135302 199958 143412 200018
rect 133183 199914 133249 199919
rect 127157 199880 128370 199882
rect 127157 199824 127162 199880
rect 127218 199824 128370 199880
rect 127157 199822 128370 199824
rect 131021 199882 131087 199885
rect 131849 199882 131915 199885
rect 131021 199880 131915 199882
rect 131021 199824 131026 199880
rect 131082 199824 131854 199880
rect 131910 199824 131915 199880
rect 131021 199822 131915 199824
rect 127157 199819 127223 199822
rect 131021 199819 131087 199822
rect 131849 199819 131915 199822
rect 132033 199882 132099 199885
rect 133183 199882 133188 199914
rect 132033 199880 133188 199882
rect 132033 199824 132038 199880
rect 132094 199858 133188 199880
rect 133244 199858 133249 199914
rect 133551 199916 133617 199919
rect 133827 199916 133893 199919
rect 133551 199914 133660 199916
rect 132094 199853 133249 199858
rect 133367 199882 133433 199885
rect 133367 199880 133476 199882
rect 132094 199824 133246 199853
rect 132033 199822 133246 199824
rect 133367 199824 133372 199880
rect 133428 199824 133476 199880
rect 133551 199858 133556 199914
rect 133612 199884 133660 199914
rect 133827 199914 133950 199916
rect 133827 199884 133832 199914
rect 133888 199884 133950 199914
rect 135115 199914 135181 199919
rect 134195 199884 134261 199885
rect 133612 199858 133644 199884
rect 133551 199853 133644 199858
rect 132033 199819 132099 199822
rect 133367 199819 133476 199824
rect 133600 199822 133644 199853
rect 133638 199820 133644 199822
rect 133708 199820 133714 199884
rect 133822 199820 133828 199884
rect 133892 199856 133950 199884
rect 134190 199882 134196 199884
rect 133892 199820 133898 199856
rect 134104 199822 134196 199882
rect 134190 199820 134196 199822
rect 134260 199820 134266 199884
rect 134379 199880 134445 199885
rect 134379 199824 134384 199880
rect 134440 199824 134445 199880
rect 134195 199819 134261 199820
rect 134379 199819 134445 199824
rect 134747 199880 134813 199885
rect 135115 199884 135120 199914
rect 135176 199884 135181 199914
rect 134747 199824 134752 199880
rect 134808 199824 134813 199880
rect 134747 199819 134813 199824
rect 135110 199820 135116 199884
rect 135180 199882 135186 199884
rect 135180 199822 135238 199882
rect 135180 199820 135186 199822
rect 126145 199746 126211 199749
rect 133416 199746 133476 199819
rect 134382 199746 134442 199819
rect 126145 199744 133476 199746
rect 126145 199688 126150 199744
rect 126206 199688 133476 199744
rect 126145 199686 133476 199688
rect 133646 199686 134442 199746
rect 126145 199683 126211 199686
rect 118693 199610 118759 199613
rect 131941 199610 132007 199613
rect 118693 199608 132007 199610
rect 118693 199552 118698 199608
rect 118754 199552 131946 199608
rect 132002 199552 132007 199608
rect 118693 199550 132007 199552
rect 118693 199547 118759 199550
rect 131941 199547 132007 199550
rect 133137 199610 133203 199613
rect 133646 199610 133706 199686
rect 133137 199608 133706 199610
rect 133137 199552 133142 199608
rect 133198 199552 133706 199608
rect 133137 199550 133706 199552
rect 134057 199610 134123 199613
rect 134750 199610 134810 199819
rect 134057 199608 134810 199610
rect 134057 199552 134062 199608
rect 134118 199552 134810 199608
rect 134057 199550 134810 199552
rect 135302 199610 135362 199958
rect 135483 199882 135549 199885
rect 135440 199880 135549 199882
rect 135440 199824 135488 199880
rect 135544 199824 135549 199880
rect 135440 199819 135549 199824
rect 135667 199882 135733 199885
rect 136214 199882 136220 199884
rect 135667 199880 136220 199882
rect 135667 199824 135672 199880
rect 135728 199824 136220 199880
rect 135667 199822 136220 199824
rect 135667 199819 135733 199822
rect 136214 199820 136220 199822
rect 136284 199820 136290 199884
rect 136495 199882 136561 199885
rect 136863 199882 136929 199885
rect 137875 199882 137941 199885
rect 136452 199880 136561 199882
rect 136452 199824 136500 199880
rect 136556 199824 136561 199880
rect 136452 199819 136561 199824
rect 136820 199880 136929 199882
rect 136820 199824 136868 199880
rect 136924 199824 136929 199880
rect 136820 199819 136929 199824
rect 137372 199880 137941 199882
rect 137372 199824 137880 199880
rect 137936 199824 137941 199880
rect 137372 199822 137941 199824
rect 135440 199749 135500 199819
rect 135437 199744 135503 199749
rect 135943 199746 136009 199749
rect 136452 199748 136512 199819
rect 135437 199688 135442 199744
rect 135498 199688 135503 199744
rect 135437 199683 135503 199688
rect 135670 199744 136009 199746
rect 135670 199688 135948 199744
rect 136004 199688 136009 199744
rect 135670 199686 136009 199688
rect 135529 199610 135595 199613
rect 135302 199608 135595 199610
rect 135302 199552 135534 199608
rect 135590 199552 135595 199608
rect 135302 199550 135595 199552
rect 135670 199610 135730 199686
rect 135943 199683 136009 199686
rect 136398 199684 136404 199748
rect 136468 199686 136512 199748
rect 136468 199684 136474 199686
rect 136820 199613 136880 199819
rect 135846 199610 135852 199612
rect 135670 199550 135852 199610
rect 133137 199547 133203 199550
rect 134057 199547 134123 199550
rect 135529 199547 135595 199550
rect 135846 199548 135852 199550
rect 135916 199548 135922 199612
rect 136817 199608 136883 199613
rect 136817 199552 136822 199608
rect 136878 199552 136883 199608
rect 136817 199547 136883 199552
rect 137372 199610 137432 199822
rect 137875 199819 137941 199822
rect 138151 199882 138217 199885
rect 138427 199884 138493 199885
rect 138151 199880 138352 199882
rect 138151 199824 138156 199880
rect 138212 199824 138352 199880
rect 138151 199822 138352 199824
rect 138151 199819 138217 199822
rect 138292 199748 138352 199822
rect 138422 199820 138428 199884
rect 138492 199882 138498 199884
rect 138492 199822 138584 199882
rect 138492 199820 138498 199822
rect 138790 199820 138796 199884
rect 138860 199882 138866 199884
rect 139071 199882 139137 199885
rect 139347 199884 139413 199885
rect 139342 199882 139348 199884
rect 138860 199880 139137 199882
rect 138860 199824 139076 199880
rect 139132 199824 139137 199880
rect 138860 199822 139137 199824
rect 139256 199822 139348 199882
rect 138860 199820 138866 199822
rect 138427 199819 138493 199820
rect 139071 199819 139137 199822
rect 139342 199820 139348 199822
rect 139412 199820 139418 199884
rect 139531 199880 139597 199885
rect 140083 199884 140149 199885
rect 140267 199884 140333 199885
rect 140078 199882 140084 199884
rect 139531 199824 139536 199880
rect 139592 199824 139597 199880
rect 139347 199819 139413 199820
rect 139531 199819 139597 199824
rect 139992 199822 140084 199882
rect 140078 199820 140084 199822
rect 140148 199820 140154 199884
rect 140262 199820 140268 199884
rect 140332 199882 140338 199884
rect 140332 199822 140424 199882
rect 140332 199820 140338 199822
rect 140998 199820 141004 199884
rect 141068 199882 141074 199884
rect 141463 199882 141529 199885
rect 141647 199882 141713 199885
rect 141068 199880 141529 199882
rect 141068 199824 141468 199880
rect 141524 199824 141529 199880
rect 141068 199822 141529 199824
rect 141068 199820 141074 199822
rect 140083 199819 140149 199820
rect 140267 199819 140333 199820
rect 141463 199819 141529 199822
rect 141604 199880 141713 199882
rect 141604 199824 141652 199880
rect 141708 199824 141713 199880
rect 141604 199819 141713 199824
rect 142107 199880 142173 199885
rect 142475 199884 142541 199885
rect 142470 199882 142476 199884
rect 142107 199824 142112 199880
rect 142168 199824 142173 199880
rect 142107 199819 142173 199824
rect 142384 199822 142476 199882
rect 142470 199820 142476 199822
rect 142540 199820 142546 199884
rect 142935 199882 143001 199885
rect 143211 199882 143277 199885
rect 143352 199882 143412 199958
rect 146431 199916 146497 199919
rect 146431 199914 146540 199916
rect 142935 199880 143044 199882
rect 142935 199824 142940 199880
rect 142996 199824 143044 199880
rect 142475 199819 142541 199820
rect 142935 199819 143044 199824
rect 143211 199880 143412 199882
rect 143211 199824 143216 199880
rect 143272 199824 143412 199880
rect 143211 199822 143412 199824
rect 144499 199882 144565 199885
rect 144678 199882 144684 199884
rect 144499 199880 144684 199882
rect 144499 199824 144504 199880
rect 144560 199824 144684 199880
rect 144499 199822 144684 199824
rect 143211 199819 143277 199822
rect 144499 199819 144565 199822
rect 144678 199820 144684 199822
rect 144748 199820 144754 199884
rect 145230 199820 145236 199884
rect 145300 199882 145306 199884
rect 145787 199882 145853 199885
rect 145300 199880 145853 199882
rect 145300 199824 145792 199880
rect 145848 199824 145853 199880
rect 146431 199858 146436 199914
rect 146492 199884 146540 199914
rect 146707 199914 146773 199919
rect 146492 199858 146524 199884
rect 146431 199853 146524 199858
rect 145300 199822 145853 199824
rect 146480 199822 146524 199853
rect 145300 199820 145306 199822
rect 145787 199819 145853 199822
rect 146518 199820 146524 199822
rect 146588 199820 146594 199884
rect 146707 199858 146712 199914
rect 146768 199858 146773 199914
rect 146707 199853 146773 199858
rect 147075 199914 147141 199919
rect 147075 199858 147080 199914
rect 147136 199858 147141 199914
rect 147075 199853 147141 199858
rect 147351 199916 147417 199919
rect 147351 199914 147460 199916
rect 147351 199858 147356 199914
rect 147412 199884 147460 199914
rect 148179 199914 148245 199919
rect 147412 199858 147444 199884
rect 147351 199853 147444 199858
rect 138238 199684 138244 199748
rect 138308 199686 138352 199748
rect 138308 199684 138314 199686
rect 138606 199684 138612 199748
rect 138676 199746 138682 199748
rect 139534 199746 139594 199819
rect 138676 199686 139594 199746
rect 138676 199684 138682 199686
rect 139710 199684 139716 199748
rect 139780 199746 139786 199748
rect 140221 199746 140287 199749
rect 139780 199744 140287 199746
rect 139780 199688 140226 199744
rect 140282 199688 140287 199744
rect 139780 199686 140287 199688
rect 139780 199684 139786 199686
rect 140221 199683 140287 199686
rect 141366 199684 141372 199748
rect 141436 199746 141442 199748
rect 141604 199746 141664 199819
rect 141436 199686 141664 199746
rect 141436 199684 141442 199686
rect 137921 199610 137987 199613
rect 137372 199608 137987 199610
rect 137372 199552 137926 199608
rect 137982 199552 137987 199608
rect 137372 199550 137987 199552
rect 137921 199547 137987 199550
rect 140037 199610 140103 199613
rect 142110 199610 142170 199819
rect 142429 199746 142495 199749
rect 140037 199608 142170 199610
rect 140037 199552 140042 199608
rect 140098 199552 142170 199608
rect 140037 199550 142170 199552
rect 142294 199744 142495 199746
rect 142294 199688 142434 199744
rect 142490 199688 142495 199744
rect 142294 199686 142495 199688
rect 142984 199748 143044 199819
rect 142984 199686 143028 199748
rect 142294 199613 142354 199686
rect 142429 199683 142495 199686
rect 143022 199684 143028 199686
rect 143092 199684 143098 199748
rect 143257 199746 143323 199749
rect 143942 199746 143948 199748
rect 143257 199744 143948 199746
rect 143257 199688 143262 199744
rect 143318 199688 143948 199744
rect 143257 199686 143948 199688
rect 143257 199683 143323 199686
rect 143942 199684 143948 199686
rect 144012 199684 144018 199748
rect 146710 199746 146770 199853
rect 147078 199749 147138 199853
rect 147400 199822 147444 199853
rect 147438 199820 147444 199822
rect 147508 199820 147514 199884
rect 147990 199820 147996 199884
rect 148060 199882 148066 199884
rect 148179 199882 148184 199914
rect 148060 199858 148184 199882
rect 148240 199858 148245 199914
rect 148060 199853 148245 199858
rect 148060 199822 148242 199853
rect 148060 199820 148066 199822
rect 146845 199746 146911 199749
rect 146710 199744 146911 199746
rect 146710 199688 146850 199744
rect 146906 199688 146911 199744
rect 146710 199686 146911 199688
rect 146845 199683 146911 199686
rect 147029 199744 147138 199749
rect 147029 199688 147034 199744
rect 147090 199688 147138 199744
rect 147029 199686 147138 199688
rect 147029 199683 147095 199686
rect 148174 199684 148180 199748
rect 148244 199746 148250 199748
rect 148731 199746 148797 199749
rect 148244 199744 148797 199746
rect 148244 199688 148736 199744
rect 148792 199688 148797 199744
rect 148244 199686 148797 199688
rect 148244 199684 148250 199686
rect 148731 199683 148797 199686
rect 142294 199608 142403 199613
rect 142294 199552 142342 199608
rect 142398 199552 142403 199608
rect 142294 199550 142403 199552
rect 140037 199547 140103 199550
rect 142337 199547 142403 199550
rect 143206 199548 143212 199612
rect 143276 199610 143282 199612
rect 143441 199610 143507 199613
rect 143276 199608 143507 199610
rect 143276 199552 143446 199608
rect 143502 199552 143507 199608
rect 143276 199550 143507 199552
rect 143276 199548 143282 199550
rect 143441 199547 143507 199550
rect 143574 199548 143580 199612
rect 143644 199610 143650 199612
rect 144729 199610 144795 199613
rect 143644 199608 144795 199610
rect 143644 199552 144734 199608
rect 144790 199552 144795 199608
rect 143644 199550 144795 199552
rect 143644 199548 143650 199550
rect 144729 199547 144795 199550
rect 146569 199610 146635 199613
rect 146886 199610 146892 199612
rect 146569 199608 146892 199610
rect 146569 199552 146574 199608
rect 146630 199552 146892 199608
rect 146569 199550 146892 199552
rect 146569 199547 146635 199550
rect 146886 199548 146892 199550
rect 146956 199548 146962 199612
rect 147305 199610 147371 199613
rect 147857 199610 147923 199613
rect 147305 199608 147923 199610
rect 147305 199552 147310 199608
rect 147366 199552 147862 199608
rect 147918 199552 147923 199608
rect 147305 199550 147923 199552
rect 148872 199610 148932 200094
rect 152322 200094 152596 200154
rect 152322 199919 152382 200094
rect 152590 200092 152596 200094
rect 152660 200092 152666 200156
rect 163446 200154 163452 200156
rect 157934 200094 163452 200154
rect 150663 199916 150729 199919
rect 151951 199916 152017 199919
rect 152135 199916 152201 199919
rect 150620 199914 150729 199916
rect 149007 199882 149073 199885
rect 149467 199884 149533 199885
rect 149462 199882 149468 199884
rect 149007 199880 149116 199882
rect 149007 199824 149012 199880
rect 149068 199824 149116 199880
rect 149007 199819 149116 199824
rect 149376 199822 149468 199882
rect 149462 199820 149468 199822
rect 149532 199820 149538 199884
rect 150014 199820 150020 199884
rect 150084 199882 150090 199884
rect 150295 199882 150361 199885
rect 150620 199884 150668 199914
rect 150084 199880 150361 199882
rect 150084 199824 150300 199880
rect 150356 199824 150361 199880
rect 150084 199822 150361 199824
rect 150084 199820 150090 199822
rect 149467 199819 149533 199820
rect 150295 199819 150361 199822
rect 150566 199820 150572 199884
rect 150636 199858 150668 199884
rect 150724 199858 150729 199914
rect 151908 199914 152017 199916
rect 150636 199853 150729 199858
rect 150636 199822 150680 199853
rect 150636 199820 150642 199822
rect 151118 199820 151124 199884
rect 151188 199882 151194 199884
rect 151908 199882 151956 199914
rect 151188 199858 151956 199882
rect 152012 199858 152017 199914
rect 151188 199853 152017 199858
rect 152092 199914 152201 199916
rect 152092 199858 152140 199914
rect 152196 199858 152201 199914
rect 152092 199853 152201 199858
rect 152319 199914 152385 199919
rect 152319 199858 152324 199914
rect 152380 199858 152385 199914
rect 152963 199914 153029 199919
rect 152687 199882 152753 199885
rect 152963 199884 152968 199914
rect 153024 199884 153029 199914
rect 153607 199916 153673 199919
rect 155815 199916 155881 199919
rect 156551 199916 156617 199919
rect 153607 199914 153946 199916
rect 152319 199853 152385 199858
rect 152506 199880 152753 199882
rect 151188 199822 151968 199853
rect 151188 199820 151194 199822
rect 149056 199749 149116 199819
rect 152092 199749 152152 199853
rect 152506 199824 152692 199880
rect 152748 199824 152753 199880
rect 152506 199822 152753 199824
rect 149053 199744 149119 199749
rect 149053 199688 149058 199744
rect 149114 199688 149119 199744
rect 149053 199683 149119 199688
rect 151491 199744 151557 199749
rect 151905 199748 151971 199749
rect 151491 199688 151496 199744
rect 151552 199688 151557 199744
rect 151491 199683 151557 199688
rect 151854 199684 151860 199748
rect 151924 199746 151971 199748
rect 151924 199744 152016 199746
rect 151966 199688 152016 199744
rect 151924 199686 152016 199688
rect 152089 199744 152155 199749
rect 152089 199688 152094 199744
rect 152150 199688 152155 199744
rect 151924 199684 151971 199686
rect 151905 199683 151971 199684
rect 152089 199683 152155 199688
rect 152222 199684 152228 199748
rect 152292 199746 152298 199748
rect 152365 199746 152431 199749
rect 152292 199744 152431 199746
rect 152292 199688 152370 199744
rect 152426 199688 152431 199744
rect 152292 199686 152431 199688
rect 152506 199746 152566 199822
rect 152687 199819 152753 199822
rect 152958 199820 152964 199884
rect 153028 199882 153034 199884
rect 153028 199822 153086 199882
rect 153607 199858 153612 199914
rect 153668 199884 153946 199914
rect 155542 199914 155881 199916
rect 153668 199858 153884 199884
rect 153607 199856 153884 199858
rect 153607 199853 153673 199856
rect 153028 199820 153034 199822
rect 153878 199820 153884 199856
rect 153948 199820 153954 199884
rect 154062 199820 154068 199884
rect 154132 199882 154138 199884
rect 154527 199882 154593 199885
rect 154132 199880 154593 199882
rect 154132 199824 154532 199880
rect 154588 199824 154593 199880
rect 154132 199822 154593 199824
rect 154132 199820 154138 199822
rect 154527 199819 154593 199822
rect 155542 199858 155820 199914
rect 155876 199858 155881 199914
rect 155542 199856 155881 199858
rect 152641 199746 152707 199749
rect 153929 199746 153995 199749
rect 152506 199744 152707 199746
rect 152506 199688 152646 199744
rect 152702 199688 152707 199744
rect 152506 199686 152707 199688
rect 152292 199684 152298 199686
rect 152365 199683 152431 199686
rect 152641 199683 152707 199686
rect 152782 199744 153995 199746
rect 152782 199688 153934 199744
rect 153990 199688 153995 199744
rect 152782 199686 153995 199688
rect 155542 199746 155602 199856
rect 155815 199853 155881 199856
rect 156416 199914 156617 199916
rect 156416 199858 156556 199914
rect 156612 199858 156617 199914
rect 157195 199914 157261 199919
rect 157011 199884 157077 199885
rect 157006 199882 157012 199884
rect 156416 199856 156617 199858
rect 155769 199746 155835 199749
rect 155542 199744 155835 199746
rect 155542 199688 155774 199744
rect 155830 199688 155835 199744
rect 155542 199686 155835 199688
rect 156416 199746 156476 199856
rect 156551 199853 156617 199856
rect 156920 199822 157012 199882
rect 157006 199820 157012 199822
rect 157076 199820 157082 199884
rect 157195 199858 157200 199914
rect 157256 199882 157261 199914
rect 157374 199882 157380 199884
rect 157256 199858 157380 199882
rect 157195 199853 157380 199858
rect 157198 199822 157380 199853
rect 157374 199820 157380 199822
rect 157444 199820 157450 199884
rect 157011 199819 157077 199820
rect 157934 199749 157994 200094
rect 163446 200092 163452 200094
rect 163516 200092 163522 200156
rect 164190 200094 170368 200154
rect 161798 199958 162916 200018
rect 158299 199914 158365 199919
rect 158943 199916 159009 199919
rect 158299 199884 158304 199914
rect 158360 199884 158365 199914
rect 158670 199914 159009 199916
rect 158294 199820 158300 199884
rect 158364 199882 158370 199884
rect 158364 199822 158422 199882
rect 158670 199858 158948 199914
rect 159004 199858 159009 199914
rect 158670 199856 159009 199858
rect 158364 199820 158370 199822
rect 156597 199746 156663 199749
rect 156416 199744 156663 199746
rect 156416 199688 156602 199744
rect 156658 199688 156663 199744
rect 156416 199686 156663 199688
rect 151494 199613 151554 199683
rect 150249 199610 150315 199613
rect 148872 199608 150315 199610
rect 148872 199552 150254 199608
rect 150310 199552 150315 199608
rect 148872 199550 150315 199552
rect 147305 199547 147371 199550
rect 147857 199547 147923 199550
rect 150249 199547 150315 199550
rect 150709 199610 150775 199613
rect 151302 199610 151308 199612
rect 150709 199608 151308 199610
rect 150709 199552 150714 199608
rect 150770 199552 151308 199608
rect 150709 199550 151308 199552
rect 150709 199547 150775 199550
rect 151302 199548 151308 199550
rect 151372 199548 151378 199612
rect 151445 199608 151554 199613
rect 151445 199552 151450 199608
rect 151506 199552 151554 199608
rect 151445 199550 151554 199552
rect 151629 199610 151695 199613
rect 152782 199610 152842 199686
rect 153929 199683 153995 199686
rect 155769 199683 155835 199686
rect 156597 199683 156663 199686
rect 156781 199748 156847 199749
rect 156781 199744 156828 199748
rect 156892 199746 156898 199748
rect 156781 199688 156786 199744
rect 156781 199684 156828 199688
rect 156892 199686 156938 199746
rect 157885 199744 157994 199749
rect 157885 199688 157890 199744
rect 157946 199688 157994 199744
rect 157885 199686 157994 199688
rect 156892 199684 156898 199686
rect 156781 199683 156847 199684
rect 157885 199683 157951 199686
rect 158110 199684 158116 199748
rect 158180 199746 158186 199748
rect 158529 199746 158595 199749
rect 158180 199744 158595 199746
rect 158180 199688 158534 199744
rect 158590 199688 158595 199744
rect 158180 199686 158595 199688
rect 158180 199684 158186 199686
rect 158529 199683 158595 199686
rect 151629 199608 152842 199610
rect 151629 199552 151634 199608
rect 151690 199552 152842 199608
rect 151629 199550 152842 199552
rect 152917 199612 152983 199613
rect 153377 199612 153443 199613
rect 152917 199608 152964 199612
rect 153028 199610 153034 199612
rect 153326 199610 153332 199612
rect 152917 199552 152922 199608
rect 151445 199547 151511 199550
rect 151629 199547 151695 199550
rect 152917 199548 152964 199552
rect 153028 199550 153074 199610
rect 153286 199550 153332 199610
rect 153396 199608 153443 199612
rect 153438 199552 153443 199608
rect 153028 199548 153034 199550
rect 153326 199548 153332 199550
rect 153396 199548 153443 199552
rect 154246 199548 154252 199612
rect 154316 199610 154322 199612
rect 154389 199610 154455 199613
rect 154316 199608 154455 199610
rect 154316 199552 154394 199608
rect 154450 199552 154455 199608
rect 154316 199550 154455 199552
rect 154316 199548 154322 199550
rect 152917 199547 152983 199548
rect 153377 199547 153443 199548
rect 154389 199547 154455 199550
rect 156638 199548 156644 199612
rect 156708 199610 156714 199612
rect 157149 199610 157215 199613
rect 156708 199608 157215 199610
rect 156708 199552 157154 199608
rect 157210 199552 157215 199608
rect 156708 199550 157215 199552
rect 156708 199548 156714 199550
rect 157149 199547 157215 199550
rect 158253 199610 158319 199613
rect 158670 199610 158730 199856
rect 158943 199853 159009 199856
rect 159219 199914 159285 199919
rect 159219 199858 159224 199914
rect 159280 199858 159285 199914
rect 160231 199916 160297 199919
rect 160599 199916 160665 199919
rect 160231 199914 160340 199916
rect 159219 199853 159285 199858
rect 158253 199608 158730 199610
rect 158253 199552 158258 199608
rect 158314 199552 158730 199608
rect 158253 199550 158730 199552
rect 159222 199613 159282 199853
rect 159398 199820 159404 199884
rect 159468 199882 159474 199884
rect 159955 199882 160021 199885
rect 159468 199880 160021 199882
rect 159468 199824 159960 199880
rect 160016 199824 160021 199880
rect 160231 199858 160236 199914
rect 160292 199884 160340 199914
rect 160556 199914 160665 199916
rect 160292 199858 160324 199884
rect 160231 199853 160324 199858
rect 159468 199822 160021 199824
rect 160280 199822 160324 199853
rect 159468 199820 159474 199822
rect 159955 199819 160021 199822
rect 160318 199820 160324 199822
rect 160388 199820 160394 199884
rect 160556 199858 160604 199914
rect 160660 199858 160665 199914
rect 160556 199853 160665 199858
rect 161243 199914 161309 199919
rect 161243 199858 161248 199914
rect 161304 199858 161309 199914
rect 161243 199853 161309 199858
rect 160556 199749 160616 199853
rect 159449 199746 159515 199749
rect 159582 199746 159588 199748
rect 159449 199744 159588 199746
rect 159449 199688 159454 199744
rect 159510 199688 159588 199744
rect 159449 199686 159588 199688
rect 159449 199683 159515 199686
rect 159582 199684 159588 199686
rect 159652 199684 159658 199748
rect 160553 199744 160619 199749
rect 160553 199688 160558 199744
rect 160614 199688 160619 199744
rect 160553 199683 160619 199688
rect 161246 199746 161306 199853
rect 161473 199746 161539 199749
rect 161246 199744 161539 199746
rect 161246 199688 161478 199744
rect 161534 199688 161539 199744
rect 161246 199686 161539 199688
rect 161473 199683 161539 199686
rect 161657 199746 161723 199749
rect 161798 199746 161858 199958
rect 161974 199820 161980 199884
rect 162044 199882 162050 199884
rect 162623 199882 162689 199885
rect 162044 199880 162689 199882
rect 162044 199824 162628 199880
rect 162684 199824 162689 199880
rect 162044 199822 162689 199824
rect 162856 199882 162916 199958
rect 163262 199956 163268 200020
rect 163332 200018 163338 200020
rect 164190 200018 164250 200094
rect 166574 200018 166580 200020
rect 163332 199958 164250 200018
rect 165892 199958 166580 200018
rect 163332 199956 163338 199958
rect 165199 199916 165265 199919
rect 165156 199914 165265 199916
rect 163543 199882 163609 199885
rect 164003 199884 164069 199885
rect 163998 199882 164004 199884
rect 162856 199880 163609 199882
rect 162856 199824 163548 199880
rect 163604 199824 163609 199880
rect 162856 199822 163609 199824
rect 163912 199822 164004 199882
rect 162044 199820 162050 199822
rect 162623 199819 162689 199822
rect 163543 199819 163609 199822
rect 163998 199820 164004 199822
rect 164068 199820 164074 199884
rect 164550 199820 164556 199884
rect 164620 199882 164626 199884
rect 165156 199882 165204 199914
rect 164620 199858 165204 199882
rect 165260 199858 165265 199914
rect 164620 199853 165265 199858
rect 165659 199882 165725 199885
rect 165892 199882 165952 199958
rect 166574 199956 166580 199958
rect 166644 199956 166650 200020
rect 166855 199916 166921 199919
rect 166855 199914 167102 199916
rect 165659 199880 165952 199882
rect 164620 199822 165216 199853
rect 165659 199824 165664 199880
rect 165720 199824 165952 199880
rect 165659 199822 165952 199824
rect 166027 199880 166093 199885
rect 166027 199824 166032 199880
rect 166088 199824 166093 199880
rect 164620 199820 164626 199822
rect 164003 199819 164069 199820
rect 165659 199819 165725 199822
rect 166027 199819 166093 199824
rect 166211 199882 166277 199885
rect 166390 199882 166396 199884
rect 166211 199880 166396 199882
rect 166211 199824 166216 199880
rect 166272 199824 166396 199880
rect 166211 199822 166396 199824
rect 166211 199819 166277 199822
rect 166390 199820 166396 199822
rect 166460 199820 166466 199884
rect 166579 199880 166645 199885
rect 166579 199824 166584 199880
rect 166640 199824 166645 199880
rect 166855 199858 166860 199914
rect 166916 199858 167102 199914
rect 167315 199914 167381 199919
rect 167315 199884 167320 199914
rect 167376 199884 167381 199914
rect 167499 199914 167565 199919
rect 166855 199856 167102 199858
rect 166855 199853 166921 199856
rect 166579 199819 166645 199824
rect 161657 199744 161858 199746
rect 161657 199688 161662 199744
rect 161718 199688 161858 199744
rect 161657 199686 161858 199688
rect 161657 199683 161723 199686
rect 162526 199684 162532 199748
rect 162596 199746 162602 199748
rect 165153 199746 165219 199749
rect 166030 199748 166090 199819
rect 162596 199744 165219 199746
rect 162596 199688 165158 199744
rect 165214 199688 165219 199744
rect 162596 199686 165219 199688
rect 162596 199684 162602 199686
rect 165153 199683 165219 199686
rect 166022 199684 166028 199748
rect 166092 199684 166098 199748
rect 166206 199684 166212 199748
rect 166276 199746 166282 199748
rect 166582 199746 166642 199819
rect 166276 199686 166642 199746
rect 166809 199746 166875 199749
rect 167042 199746 167102 199856
rect 167310 199820 167316 199884
rect 167380 199882 167386 199884
rect 167380 199822 167438 199882
rect 167499 199858 167504 199914
rect 167560 199858 167565 199914
rect 169891 199914 169957 199919
rect 168603 199884 168669 199885
rect 167499 199853 167565 199858
rect 167380 199820 167386 199822
rect 167502 199749 167562 199853
rect 168598 199820 168604 199884
rect 168668 199882 168674 199884
rect 168668 199822 168760 199882
rect 168668 199820 168674 199822
rect 168966 199820 168972 199884
rect 169036 199882 169042 199884
rect 169247 199882 169313 199885
rect 169036 199880 169313 199882
rect 169036 199824 169252 199880
rect 169308 199824 169313 199880
rect 169036 199822 169313 199824
rect 169036 199820 169042 199822
rect 168603 199819 168669 199820
rect 169247 199819 169313 199822
rect 169431 199882 169497 199885
rect 169431 199880 169770 199882
rect 169431 199824 169436 199880
rect 169492 199824 169770 199880
rect 169891 199858 169896 199914
rect 169952 199858 169957 199914
rect 169891 199853 169957 199858
rect 169431 199822 169770 199824
rect 169431 199819 169497 199822
rect 166809 199744 167102 199746
rect 166809 199688 166814 199744
rect 166870 199688 167102 199744
rect 166809 199686 167102 199688
rect 167453 199744 167562 199749
rect 167453 199688 167458 199744
rect 167514 199688 167562 199744
rect 167453 199686 167562 199688
rect 166276 199684 166282 199686
rect 166809 199683 166875 199686
rect 167453 199683 167519 199686
rect 169334 199684 169340 199748
rect 169404 199746 169410 199748
rect 169710 199746 169770 199822
rect 169894 199749 169954 199853
rect 169404 199686 169770 199746
rect 169845 199744 169954 199749
rect 169845 199688 169850 199744
rect 169906 199688 169954 199744
rect 169845 199686 169954 199688
rect 169404 199684 169410 199686
rect 169845 199683 169911 199686
rect 170308 199613 170368 200094
rect 170990 200092 170996 200156
rect 171060 200154 171066 200156
rect 180517 200154 180583 200157
rect 209814 200154 209820 200156
rect 171060 200094 172530 200154
rect 171060 200092 171066 200094
rect 172470 199919 172530 200094
rect 173896 200094 175474 200154
rect 173198 199956 173204 200020
rect 173268 200018 173274 200020
rect 173268 199956 173312 200018
rect 170627 199914 170693 199919
rect 170627 199884 170632 199914
rect 170688 199884 170693 199914
rect 170903 199916 170969 199919
rect 171639 199916 171705 199919
rect 170903 199914 171012 199916
rect 170622 199820 170628 199884
rect 170692 199882 170698 199884
rect 170692 199822 170750 199882
rect 170903 199858 170908 199914
rect 170964 199882 171012 199914
rect 171596 199914 171705 199916
rect 171358 199882 171364 199884
rect 170964 199858 171364 199882
rect 170903 199853 171364 199858
rect 170952 199822 171364 199853
rect 170692 199820 170698 199822
rect 171358 199820 171364 199822
rect 171428 199820 171434 199884
rect 171596 199858 171644 199914
rect 171700 199858 171705 199914
rect 171596 199853 171705 199858
rect 172007 199916 172073 199919
rect 172007 199914 172208 199916
rect 172007 199858 172012 199914
rect 172068 199882 172208 199914
rect 172467 199914 172533 199919
rect 172278 199882 172284 199884
rect 172068 199858 172284 199882
rect 172007 199856 172284 199858
rect 172007 199853 172073 199856
rect 171317 199746 171383 199749
rect 171596 199746 171656 199853
rect 172148 199822 172284 199856
rect 172278 199820 172284 199822
rect 172348 199820 172354 199884
rect 172467 199858 172472 199914
rect 172528 199858 172533 199914
rect 172467 199853 172533 199858
rect 172743 199882 172809 199885
rect 173111 199882 173177 199885
rect 173252 199882 173312 199956
rect 173896 199919 173956 200094
rect 172743 199880 172944 199882
rect 172743 199824 172748 199880
rect 172804 199824 172944 199880
rect 172743 199822 172944 199824
rect 172743 199819 172809 199822
rect 171317 199744 171656 199746
rect 171317 199688 171322 199744
rect 171378 199688 171656 199744
rect 171317 199686 171656 199688
rect 172884 199746 172944 199822
rect 173111 199880 173312 199882
rect 173111 199824 173116 199880
rect 173172 199824 173312 199880
rect 173847 199914 173956 199919
rect 173847 199858 173852 199914
rect 173908 199858 173956 199914
rect 174307 199914 174373 199919
rect 174307 199884 174312 199914
rect 174368 199884 174373 199914
rect 174491 199914 174557 199919
rect 173847 199856 173956 199858
rect 173847 199853 173913 199856
rect 173111 199822 173312 199824
rect 173111 199819 173177 199822
rect 174302 199820 174308 199884
rect 174372 199882 174378 199884
rect 174372 199822 174430 199882
rect 174491 199858 174496 199914
rect 174552 199858 174557 199914
rect 174675 199914 174741 199919
rect 174675 199884 174680 199914
rect 174736 199884 174741 199914
rect 174491 199853 174557 199858
rect 174372 199820 174378 199822
rect 174494 199749 174554 199853
rect 174670 199820 174676 199884
rect 174740 199882 174746 199884
rect 174740 199822 174798 199882
rect 174740 199820 174746 199822
rect 173847 199746 173913 199749
rect 172884 199744 173913 199746
rect 172884 199688 173852 199744
rect 173908 199688 173913 199744
rect 172884 199686 173913 199688
rect 174494 199744 174603 199749
rect 174494 199688 174542 199744
rect 174598 199688 174603 199744
rect 174494 199686 174603 199688
rect 175414 199746 175474 200094
rect 175782 200094 178188 200154
rect 175782 199919 175842 200094
rect 178128 200021 178188 200094
rect 180517 200152 209820 200154
rect 180517 200096 180522 200152
rect 180578 200096 209820 200152
rect 180517 200094 209820 200096
rect 180517 200091 180583 200094
rect 209814 200092 209820 200094
rect 209884 200154 209890 200156
rect 210918 200154 210924 200156
rect 209884 200094 210924 200154
rect 209884 200092 209890 200094
rect 210918 200092 210924 200094
rect 210988 200092 210994 200156
rect 178125 200016 178191 200021
rect 178125 199960 178130 200016
rect 178186 199960 178191 200016
rect 178125 199955 178191 199960
rect 180057 200018 180123 200021
rect 180190 200018 180196 200020
rect 180057 200016 180196 200018
rect 180057 199960 180062 200016
rect 180118 199960 180196 200016
rect 180057 199958 180196 199960
rect 180057 199955 180123 199958
rect 180190 199956 180196 199958
rect 180260 199956 180266 200020
rect 175779 199914 175845 199919
rect 175779 199858 175784 199914
rect 175840 199858 175845 199914
rect 176607 199914 176673 199919
rect 175779 199853 175845 199858
rect 176326 199820 176332 199884
rect 176396 199882 176402 199884
rect 176607 199882 176612 199914
rect 176396 199858 176612 199882
rect 176668 199858 176673 199914
rect 176396 199853 176673 199858
rect 176883 199914 176949 199919
rect 176883 199858 176888 199914
rect 176944 199882 176949 199914
rect 177849 199882 177915 199885
rect 176944 199880 177915 199882
rect 176944 199858 177854 199880
rect 176883 199853 177854 199858
rect 176396 199822 176670 199853
rect 176886 199824 177854 199853
rect 177910 199824 177915 199880
rect 176886 199822 177915 199824
rect 176396 199820 176402 199822
rect 177849 199819 177915 199822
rect 178585 199746 178651 199749
rect 175414 199744 178651 199746
rect 175414 199688 178590 199744
rect 178646 199688 178651 199744
rect 175414 199686 178651 199688
rect 171317 199683 171383 199686
rect 173847 199683 173913 199686
rect 174537 199683 174603 199686
rect 178585 199683 178651 199686
rect 180241 199746 180307 199749
rect 188470 199746 188476 199748
rect 180241 199744 188476 199746
rect 180241 199688 180246 199744
rect 180302 199688 188476 199744
rect 180241 199686 188476 199688
rect 180241 199683 180307 199686
rect 188470 199684 188476 199686
rect 188540 199684 188546 199748
rect 159222 199608 159331 199613
rect 159222 199552 159270 199608
rect 159326 199552 159331 199608
rect 159222 199550 159331 199552
rect 158253 199547 158319 199550
rect 159265 199547 159331 199550
rect 160737 199610 160803 199613
rect 160870 199610 160876 199612
rect 160737 199608 160876 199610
rect 160737 199552 160742 199608
rect 160798 199552 160876 199608
rect 160737 199550 160876 199552
rect 160737 199547 160803 199550
rect 160870 199548 160876 199550
rect 160940 199548 160946 199612
rect 164509 199610 164575 199613
rect 164734 199610 164740 199612
rect 164509 199608 164740 199610
rect 164509 199552 164514 199608
rect 164570 199552 164740 199608
rect 164509 199550 164740 199552
rect 164509 199547 164575 199550
rect 164734 199548 164740 199550
rect 164804 199548 164810 199612
rect 164877 199610 164943 199613
rect 165102 199610 165108 199612
rect 164877 199608 165108 199610
rect 164877 199552 164882 199608
rect 164938 199552 165108 199608
rect 164877 199550 165108 199552
rect 164877 199547 164943 199550
rect 165102 199548 165108 199550
rect 165172 199548 165178 199612
rect 168649 199610 168715 199613
rect 169150 199610 169156 199612
rect 168649 199608 169156 199610
rect 168649 199552 168654 199608
rect 168710 199552 169156 199608
rect 168649 199550 169156 199552
rect 168649 199547 168715 199550
rect 169150 199548 169156 199550
rect 169220 199548 169226 199612
rect 169385 199610 169451 199613
rect 169518 199610 169524 199612
rect 169385 199608 169524 199610
rect 169385 199552 169390 199608
rect 169446 199552 169524 199608
rect 169385 199550 169524 199552
rect 169385 199547 169451 199550
rect 169518 199548 169524 199550
rect 169588 199548 169594 199612
rect 170305 199608 170371 199613
rect 170857 199612 170923 199613
rect 170806 199610 170812 199612
rect 170305 199552 170310 199608
rect 170366 199552 170371 199608
rect 170305 199547 170371 199552
rect 170766 199550 170812 199610
rect 170876 199608 170923 199612
rect 170918 199552 170923 199608
rect 170806 199548 170812 199550
rect 170876 199548 170923 199552
rect 170857 199547 170923 199548
rect 171685 199610 171751 199613
rect 178861 199610 178927 199613
rect 189717 199610 189783 199613
rect 171685 199608 189783 199610
rect 171685 199552 171690 199608
rect 171746 199552 178866 199608
rect 178922 199552 189722 199608
rect 189778 199552 189783 199608
rect 171685 199550 189783 199552
rect 171685 199547 171751 199550
rect 178861 199547 178927 199550
rect 189717 199547 189783 199550
rect 205582 199548 205588 199612
rect 205652 199610 205658 199612
rect 548609 199610 548675 199613
rect 205652 199608 548675 199610
rect 205652 199552 548614 199608
rect 548670 199552 548675 199608
rect 205652 199550 548675 199552
rect 205652 199548 205658 199550
rect 548609 199547 548675 199550
rect 31017 199474 31083 199477
rect 107510 199474 107516 199476
rect 31017 199472 107516 199474
rect 31017 199416 31022 199472
rect 31078 199416 107516 199472
rect 31017 199414 107516 199416
rect 31017 199411 31083 199414
rect 107510 199412 107516 199414
rect 107580 199412 107586 199476
rect 122414 199412 122420 199476
rect 122484 199474 122490 199476
rect 172605 199474 172671 199477
rect 122484 199472 172671 199474
rect 122484 199416 172610 199472
rect 172666 199416 172671 199472
rect 122484 199414 172671 199416
rect 122484 199412 122490 199414
rect 172605 199411 172671 199414
rect 175406 199412 175412 199476
rect 175476 199474 175482 199476
rect 176193 199474 176259 199477
rect 175476 199472 176259 199474
rect 175476 199416 176198 199472
rect 176254 199416 176259 199472
rect 175476 199414 176259 199416
rect 175476 199412 175482 199414
rect 176193 199411 176259 199414
rect 176326 199412 176332 199476
rect 176396 199474 176402 199476
rect 179321 199474 179387 199477
rect 176396 199472 179387 199474
rect 176396 199416 179326 199472
rect 179382 199416 179387 199472
rect 176396 199414 179387 199416
rect 176396 199412 176402 199414
rect 179321 199411 179387 199414
rect 180701 199474 180767 199477
rect 580533 199474 580599 199477
rect 180701 199472 580599 199474
rect 180701 199416 180706 199472
rect 180762 199416 580538 199472
rect 580594 199416 580599 199472
rect 180701 199414 580599 199416
rect 180701 199411 180767 199414
rect 580533 199411 580599 199414
rect 4153 199338 4219 199341
rect 161974 199338 161980 199340
rect 4153 199336 161980 199338
rect 4153 199280 4158 199336
rect 4214 199280 161980 199336
rect 4153 199278 161980 199280
rect 4153 199275 4219 199278
rect 161974 199276 161980 199278
rect 162044 199276 162050 199340
rect 162485 199338 162551 199341
rect 163262 199338 163268 199340
rect 162485 199336 163268 199338
rect 162485 199280 162490 199336
rect 162546 199280 163268 199336
rect 162485 199278 163268 199280
rect 162485 199275 162551 199278
rect 163262 199276 163268 199278
rect 163332 199276 163338 199340
rect 165889 199338 165955 199341
rect 168414 199338 168420 199340
rect 165889 199336 168420 199338
rect 165889 199280 165894 199336
rect 165950 199280 168420 199336
rect 165889 199278 168420 199280
rect 165889 199275 165955 199278
rect 168414 199276 168420 199278
rect 168484 199276 168490 199340
rect 170949 199338 171015 199341
rect 580349 199338 580415 199341
rect 170949 199336 580415 199338
rect 170949 199280 170954 199336
rect 171010 199280 580354 199336
rect 580410 199280 580415 199336
rect 170949 199278 580415 199280
rect 170949 199275 171015 199278
rect 580349 199275 580415 199278
rect 133597 199202 133663 199205
rect 136265 199202 136331 199205
rect 133597 199200 136331 199202
rect 133597 199144 133602 199200
rect 133658 199144 136270 199200
rect 136326 199144 136331 199200
rect 133597 199142 136331 199144
rect 133597 199139 133663 199142
rect 136265 199139 136331 199142
rect 137829 199202 137895 199205
rect 139301 199202 139367 199205
rect 140037 199204 140103 199205
rect 139710 199202 139716 199204
rect 137829 199200 139226 199202
rect 137829 199144 137834 199200
rect 137890 199144 139226 199200
rect 137829 199142 139226 199144
rect 137829 199139 137895 199142
rect 125593 199066 125659 199069
rect 139025 199066 139091 199069
rect 125593 199064 139091 199066
rect 125593 199008 125598 199064
rect 125654 199008 139030 199064
rect 139086 199008 139091 199064
rect 125593 199006 139091 199008
rect 139166 199066 139226 199142
rect 139301 199200 139716 199202
rect 139301 199144 139306 199200
rect 139362 199144 139716 199200
rect 139301 199142 139716 199144
rect 139301 199139 139367 199142
rect 139710 199140 139716 199142
rect 139780 199140 139786 199204
rect 140037 199202 140084 199204
rect 139992 199200 140084 199202
rect 139992 199144 140042 199200
rect 139992 199142 140084 199144
rect 140037 199140 140084 199142
rect 140148 199140 140154 199204
rect 140446 199140 140452 199204
rect 140516 199202 140522 199204
rect 144085 199202 144151 199205
rect 140516 199200 144151 199202
rect 140516 199144 144090 199200
rect 144146 199144 144151 199200
rect 140516 199142 144151 199144
rect 140516 199140 140522 199142
rect 140037 199139 140103 199140
rect 144085 199139 144151 199142
rect 150249 199202 150315 199205
rect 152641 199202 152707 199205
rect 150249 199200 152707 199202
rect 150249 199144 150254 199200
rect 150310 199144 152646 199200
rect 152702 199144 152707 199200
rect 150249 199142 152707 199144
rect 150249 199139 150315 199142
rect 152641 199139 152707 199142
rect 153101 199202 153167 199205
rect 153694 199202 153700 199204
rect 153101 199200 153700 199202
rect 153101 199144 153106 199200
rect 153162 199144 153700 199200
rect 153101 199142 153700 199144
rect 153101 199139 153167 199142
rect 153694 199140 153700 199142
rect 153764 199140 153770 199204
rect 153929 199202 153995 199205
rect 184974 199202 184980 199204
rect 153929 199200 184980 199202
rect 153929 199144 153934 199200
rect 153990 199144 184980 199200
rect 153929 199142 184980 199144
rect 153929 199139 153995 199142
rect 184974 199140 184980 199142
rect 185044 199140 185050 199204
rect 143073 199066 143139 199069
rect 139166 199064 143139 199066
rect 139166 199008 143078 199064
rect 143134 199008 143139 199064
rect 139166 199006 143139 199008
rect 125593 199003 125659 199006
rect 139025 199003 139091 199006
rect 143073 199003 143139 199006
rect 143390 199004 143396 199068
rect 143460 199066 143466 199068
rect 144729 199066 144795 199069
rect 143460 199064 144795 199066
rect 143460 199008 144734 199064
rect 144790 199008 144795 199064
rect 143460 199006 144795 199008
rect 143460 199004 143466 199006
rect 144729 199003 144795 199006
rect 150566 199004 150572 199068
rect 150636 199066 150642 199068
rect 150709 199066 150775 199069
rect 150636 199064 150775 199066
rect 150636 199008 150714 199064
rect 150770 199008 150775 199064
rect 150636 199006 150775 199008
rect 150636 199004 150642 199006
rect 150709 199003 150775 199006
rect 150985 199066 151051 199069
rect 151629 199068 151695 199069
rect 151486 199066 151492 199068
rect 150985 199064 151492 199066
rect 150985 199008 150990 199064
rect 151046 199008 151492 199064
rect 150985 199006 151492 199008
rect 150985 199003 151051 199006
rect 151486 199004 151492 199006
rect 151556 199004 151562 199068
rect 151629 199064 151676 199068
rect 151740 199066 151746 199068
rect 152089 199066 152155 199069
rect 171685 199066 171751 199069
rect 179597 199066 179663 199069
rect 180701 199066 180767 199069
rect 151629 199008 151634 199064
rect 151629 199004 151676 199008
rect 151740 199006 151786 199066
rect 152089 199064 171751 199066
rect 152089 199008 152094 199064
rect 152150 199008 171690 199064
rect 171746 199008 171751 199064
rect 152089 199006 171751 199008
rect 151740 199004 151746 199006
rect 151629 199003 151695 199004
rect 152089 199003 152155 199006
rect 171685 199003 171751 199006
rect 171918 199064 180767 199066
rect 171918 199008 179602 199064
rect 179658 199008 180706 199064
rect 180762 199008 180767 199064
rect 171918 199006 180767 199008
rect 117037 198930 117103 198933
rect 151118 198930 151124 198932
rect 117037 198928 151124 198930
rect 117037 198872 117042 198928
rect 117098 198872 151124 198928
rect 117037 198870 151124 198872
rect 117037 198867 117103 198870
rect 151118 198868 151124 198870
rect 151188 198868 151194 198932
rect 151302 198868 151308 198932
rect 151372 198930 151378 198932
rect 151629 198930 151695 198933
rect 151372 198928 151695 198930
rect 151372 198872 151634 198928
rect 151690 198872 151695 198928
rect 151372 198870 151695 198872
rect 151372 198868 151378 198870
rect 151629 198867 151695 198870
rect 151813 198930 151879 198933
rect 152038 198930 152044 198932
rect 151813 198928 152044 198930
rect 151813 198872 151818 198928
rect 151874 198872 152044 198928
rect 151813 198870 152044 198872
rect 151813 198867 151879 198870
rect 152038 198868 152044 198870
rect 152108 198868 152114 198932
rect 152273 198930 152339 198933
rect 152733 198930 152799 198933
rect 152273 198928 152799 198930
rect 152273 198872 152278 198928
rect 152334 198872 152738 198928
rect 152794 198872 152799 198928
rect 152273 198870 152799 198872
rect 152273 198867 152339 198870
rect 152733 198867 152799 198870
rect 153745 198930 153811 198933
rect 153878 198930 153884 198932
rect 153745 198928 153884 198930
rect 153745 198872 153750 198928
rect 153806 198872 153884 198928
rect 153745 198870 153884 198872
rect 153745 198867 153811 198870
rect 153878 198868 153884 198870
rect 153948 198868 153954 198932
rect 158161 198930 158227 198933
rect 158294 198930 158300 198932
rect 158161 198928 158300 198930
rect 158161 198872 158166 198928
rect 158222 198872 158300 198928
rect 158161 198870 158300 198872
rect 158161 198867 158227 198870
rect 158294 198868 158300 198870
rect 158364 198868 158370 198932
rect 164049 198930 164115 198933
rect 164877 198930 164943 198933
rect 164049 198928 164943 198930
rect 164049 198872 164054 198928
rect 164110 198872 164882 198928
rect 164938 198872 164943 198928
rect 164049 198870 164943 198872
rect 164049 198867 164115 198870
rect 164877 198867 164943 198870
rect 167637 198930 167703 198933
rect 167862 198930 167868 198932
rect 167637 198928 167868 198930
rect 167637 198872 167642 198928
rect 167698 198872 167868 198928
rect 167637 198870 167868 198872
rect 167637 198867 167703 198870
rect 167862 198868 167868 198870
rect 167932 198868 167938 198932
rect 168373 198930 168439 198933
rect 171918 198930 171978 199006
rect 179597 199003 179663 199006
rect 180701 199003 180767 199006
rect 168373 198928 171978 198930
rect 168373 198872 168378 198928
rect 168434 198872 171978 198928
rect 168373 198870 171978 198872
rect 172329 198930 172395 198933
rect 173566 198930 173572 198932
rect 172329 198928 173572 198930
rect 172329 198872 172334 198928
rect 172390 198872 173572 198928
rect 172329 198870 173572 198872
rect 168373 198867 168439 198870
rect 172329 198867 172395 198870
rect 173566 198868 173572 198870
rect 173636 198868 173642 198932
rect 178677 198930 178743 198933
rect 205582 198930 205588 198932
rect 178677 198928 205588 198930
rect 178677 198872 178682 198928
rect 178738 198872 205588 198928
rect 178677 198870 205588 198872
rect 178677 198867 178743 198870
rect 205582 198868 205588 198870
rect 205652 198930 205658 198932
rect 206134 198930 206140 198932
rect 205652 198870 206140 198930
rect 205652 198868 205658 198870
rect 206134 198868 206140 198870
rect 206204 198868 206210 198932
rect 107510 198732 107516 198796
rect 107580 198794 107586 198796
rect 135897 198794 135963 198797
rect 107580 198792 135963 198794
rect 107580 198736 135902 198792
rect 135958 198736 135963 198792
rect 107580 198734 135963 198736
rect 107580 198732 107586 198734
rect 135897 198731 135963 198734
rect 141417 198794 141483 198797
rect 142705 198794 142771 198797
rect 141417 198792 142771 198794
rect 141417 198736 141422 198792
rect 141478 198736 142710 198792
rect 142766 198736 142771 198792
rect 141417 198734 142771 198736
rect 141417 198731 141483 198734
rect 142705 198731 142771 198734
rect 142981 198794 143047 198797
rect 157885 198794 157951 198797
rect 142981 198792 157951 198794
rect 142981 198736 142986 198792
rect 143042 198736 157890 198792
rect 157946 198736 157951 198792
rect 142981 198734 157951 198736
rect 142981 198731 143047 198734
rect 157885 198731 157951 198734
rect 164734 198732 164740 198796
rect 164804 198794 164810 198796
rect 165153 198794 165219 198797
rect 164804 198792 165219 198794
rect 164804 198736 165158 198792
rect 165214 198736 165219 198792
rect 164804 198734 165219 198736
rect 164804 198732 164810 198734
rect 165153 198731 165219 198734
rect 165429 198794 165495 198797
rect 170949 198794 171015 198797
rect 177665 198794 177731 198797
rect 165429 198792 171015 198794
rect 165429 198736 165434 198792
rect 165490 198736 170954 198792
rect 171010 198736 171015 198792
rect 165429 198734 171015 198736
rect 165429 198731 165495 198734
rect 170949 198731 171015 198734
rect 172470 198792 177731 198794
rect 172470 198736 177670 198792
rect 177726 198736 177731 198792
rect 172470 198734 177731 198736
rect 137093 198658 137159 198661
rect 138790 198658 138796 198660
rect 137093 198656 138796 198658
rect 137093 198600 137098 198656
rect 137154 198600 138796 198656
rect 137093 198598 138796 198600
rect 137093 198595 137159 198598
rect 138790 198596 138796 198598
rect 138860 198596 138866 198660
rect 161933 198658 161999 198661
rect 162710 198658 162716 198660
rect 161933 198656 162716 198658
rect 161933 198600 161938 198656
rect 161994 198600 162716 198656
rect 161933 198598 162716 198600
rect 161933 198595 161999 198598
rect 162710 198596 162716 198598
rect 162780 198596 162786 198660
rect 164785 198658 164851 198661
rect 172470 198658 172530 198734
rect 177665 198731 177731 198734
rect 164785 198656 172530 198658
rect 164785 198600 164790 198656
rect 164846 198600 172530 198656
rect 164785 198598 172530 198600
rect 173249 198658 173315 198661
rect 173709 198660 173775 198661
rect 174629 198660 174695 198661
rect 173382 198658 173388 198660
rect 173249 198656 173388 198658
rect 173249 198600 173254 198656
rect 173310 198600 173388 198656
rect 173249 198598 173388 198600
rect 164785 198595 164851 198598
rect 173249 198595 173315 198598
rect 173382 198596 173388 198598
rect 173452 198596 173458 198660
rect 173709 198656 173756 198660
rect 173820 198658 173826 198660
rect 174629 198658 174676 198660
rect 173709 198600 173714 198656
rect 173709 198596 173756 198600
rect 173820 198598 173866 198658
rect 174584 198656 174676 198658
rect 174584 198600 174634 198656
rect 174584 198598 174676 198600
rect 173820 198596 173826 198598
rect 174629 198596 174676 198598
rect 174740 198596 174746 198660
rect 173709 198595 173775 198596
rect 174629 198595 174695 198596
rect 127709 198522 127775 198525
rect 137185 198522 137251 198525
rect 127709 198520 137251 198522
rect 127709 198464 127714 198520
rect 127770 198464 137190 198520
rect 137246 198464 137251 198520
rect 127709 198462 137251 198464
rect 127709 198459 127775 198462
rect 137185 198459 137251 198462
rect 138013 198522 138079 198525
rect 142245 198524 142311 198525
rect 140262 198522 140268 198524
rect 138013 198520 140268 198522
rect 138013 198464 138018 198520
rect 138074 198464 140268 198520
rect 138013 198462 140268 198464
rect 138013 198459 138079 198462
rect 140262 198460 140268 198462
rect 140332 198460 140338 198524
rect 142245 198522 142292 198524
rect 142200 198520 142292 198522
rect 142200 198464 142250 198520
rect 142200 198462 142292 198464
rect 142245 198460 142292 198462
rect 142356 198460 142362 198524
rect 144494 198460 144500 198524
rect 144564 198522 144570 198524
rect 147305 198522 147371 198525
rect 144564 198520 147371 198522
rect 144564 198464 147310 198520
rect 147366 198464 147371 198520
rect 144564 198462 147371 198464
rect 144564 198460 144570 198462
rect 142245 198459 142311 198460
rect 147305 198459 147371 198462
rect 150985 198522 151051 198525
rect 159725 198522 159791 198525
rect 150985 198520 159791 198522
rect 150985 198464 150990 198520
rect 151046 198464 159730 198520
rect 159786 198464 159791 198520
rect 150985 198462 159791 198464
rect 150985 198459 151051 198462
rect 159725 198459 159791 198462
rect 164325 198522 164391 198525
rect 180057 198522 180123 198525
rect 164325 198520 180123 198522
rect 164325 198464 164330 198520
rect 164386 198464 180062 198520
rect 180118 198464 180123 198520
rect 164325 198462 180123 198464
rect 164325 198459 164391 198462
rect 180057 198459 180123 198462
rect 133505 198386 133571 198389
rect 142153 198386 142219 198389
rect 133505 198384 142219 198386
rect 133505 198328 133510 198384
rect 133566 198328 142158 198384
rect 142214 198328 142219 198384
rect 133505 198326 142219 198328
rect 133505 198323 133571 198326
rect 142153 198323 142219 198326
rect 147070 198324 147076 198388
rect 147140 198386 147146 198388
rect 147397 198386 147463 198389
rect 147140 198384 147463 198386
rect 147140 198328 147402 198384
rect 147458 198328 147463 198384
rect 147140 198326 147463 198328
rect 147140 198324 147146 198326
rect 147397 198323 147463 198326
rect 160921 198386 160987 198389
rect 165470 198386 165476 198388
rect 160921 198384 165476 198386
rect 160921 198328 160926 198384
rect 160982 198328 165476 198384
rect 160921 198326 165476 198328
rect 160921 198323 160987 198326
rect 165470 198324 165476 198326
rect 165540 198324 165546 198388
rect 167085 198386 167151 198389
rect 180241 198386 180307 198389
rect 167085 198384 180307 198386
rect 167085 198328 167090 198384
rect 167146 198328 180246 198384
rect 180302 198328 180307 198384
rect 167085 198326 180307 198328
rect 167085 198323 167151 198326
rect 180241 198323 180307 198326
rect 124121 198250 124187 198253
rect 134609 198250 134675 198253
rect 124121 198248 134675 198250
rect 124121 198192 124126 198248
rect 124182 198192 134614 198248
rect 134670 198192 134675 198248
rect 124121 198190 134675 198192
rect 124121 198187 124187 198190
rect 134609 198187 134675 198190
rect 136633 198250 136699 198253
rect 138289 198250 138355 198253
rect 136633 198248 138355 198250
rect 136633 198192 136638 198248
rect 136694 198192 138294 198248
rect 138350 198192 138355 198248
rect 136633 198190 138355 198192
rect 136633 198187 136699 198190
rect 138289 198187 138355 198190
rect 138749 198250 138815 198253
rect 138974 198250 138980 198252
rect 138749 198248 138980 198250
rect 138749 198192 138754 198248
rect 138810 198192 138980 198248
rect 138749 198190 138980 198192
rect 138749 198187 138815 198190
rect 138974 198188 138980 198190
rect 139044 198188 139050 198252
rect 140957 198250 141023 198253
rect 141366 198250 141372 198252
rect 140957 198248 141372 198250
rect 140957 198192 140962 198248
rect 141018 198192 141372 198248
rect 140957 198190 141372 198192
rect 140957 198187 141023 198190
rect 141366 198188 141372 198190
rect 141436 198188 141442 198252
rect 159582 198188 159588 198252
rect 159652 198250 159658 198252
rect 159817 198250 159883 198253
rect 159652 198248 159883 198250
rect 159652 198192 159822 198248
rect 159878 198192 159883 198248
rect 159652 198190 159883 198192
rect 159652 198188 159658 198190
rect 159817 198187 159883 198190
rect 126881 198114 126947 198117
rect 139669 198114 139735 198117
rect 151077 198114 151143 198117
rect 126881 198112 139735 198114
rect 126881 198056 126886 198112
rect 126942 198056 139674 198112
rect 139730 198056 139735 198112
rect 126881 198054 139735 198056
rect 126881 198051 126947 198054
rect 139669 198051 139735 198054
rect 144870 198112 151143 198114
rect 144870 198056 151082 198112
rect 151138 198056 151143 198112
rect 144870 198054 151143 198056
rect 131757 197978 131823 197981
rect 135253 197978 135319 197981
rect 144870 197978 144930 198054
rect 151077 198051 151143 198054
rect 158713 198114 158779 198117
rect 158713 198112 165722 198114
rect 158713 198056 158718 198112
rect 158774 198056 165722 198112
rect 158713 198054 165722 198056
rect 158713 198051 158779 198054
rect 131757 197976 135319 197978
rect 131757 197920 131762 197976
rect 131818 197920 135258 197976
rect 135314 197920 135319 197976
rect 131757 197918 135319 197920
rect 131757 197915 131823 197918
rect 135253 197915 135319 197918
rect 137510 197918 144930 197978
rect 134374 197780 134380 197844
rect 134444 197842 134450 197844
rect 136633 197842 136699 197845
rect 134444 197840 136699 197842
rect 134444 197784 136638 197840
rect 136694 197784 136699 197840
rect 134444 197782 136699 197784
rect 134444 197780 134450 197782
rect 136633 197779 136699 197782
rect 136817 197842 136883 197845
rect 137510 197842 137570 197918
rect 147990 197916 147996 197980
rect 148060 197978 148066 197980
rect 148685 197978 148751 197981
rect 148961 197980 149027 197981
rect 148910 197978 148916 197980
rect 148060 197976 148751 197978
rect 148060 197920 148690 197976
rect 148746 197920 148751 197976
rect 148060 197918 148751 197920
rect 148870 197918 148916 197978
rect 148980 197976 149027 197980
rect 149022 197920 149027 197976
rect 148060 197916 148066 197918
rect 148685 197915 148751 197918
rect 148910 197916 148916 197918
rect 148980 197916 149027 197920
rect 148961 197915 149027 197916
rect 163221 197978 163287 197981
rect 163630 197978 163636 197980
rect 163221 197976 163636 197978
rect 163221 197920 163226 197976
rect 163282 197920 163636 197976
rect 163221 197918 163636 197920
rect 163221 197915 163287 197918
rect 163630 197916 163636 197918
rect 163700 197916 163706 197980
rect 164233 197978 164299 197981
rect 165429 197978 165495 197981
rect 164233 197976 165495 197978
rect 164233 197920 164238 197976
rect 164294 197920 165434 197976
rect 165490 197920 165495 197976
rect 164233 197918 165495 197920
rect 165662 197978 165722 198054
rect 179413 197978 179479 197981
rect 165662 197976 179479 197978
rect 165662 197920 179418 197976
rect 179474 197920 179479 197976
rect 165662 197918 179479 197920
rect 164233 197915 164299 197918
rect 165429 197915 165495 197918
rect 179413 197915 179479 197918
rect 183553 197978 183619 197981
rect 185342 197978 185348 197980
rect 183553 197976 185348 197978
rect 183553 197920 183558 197976
rect 183614 197920 185348 197976
rect 183553 197918 185348 197920
rect 183553 197915 183619 197918
rect 185342 197916 185348 197918
rect 185412 197978 185418 197980
rect 197353 197978 197419 197981
rect 185412 197976 197419 197978
rect 185412 197920 197358 197976
rect 197414 197920 197419 197976
rect 185412 197918 197419 197920
rect 185412 197916 185418 197918
rect 197353 197915 197419 197918
rect 580165 197978 580231 197981
rect 583520 197978 584960 198068
rect 580165 197976 584960 197978
rect 580165 197920 580170 197976
rect 580226 197920 584960 197976
rect 580165 197918 584960 197920
rect 580165 197915 580231 197918
rect 136817 197840 137570 197842
rect 136817 197784 136822 197840
rect 136878 197784 137570 197840
rect 136817 197782 137570 197784
rect 140865 197842 140931 197845
rect 140998 197842 141004 197844
rect 140865 197840 141004 197842
rect 140865 197784 140870 197840
rect 140926 197784 141004 197840
rect 140865 197782 141004 197784
rect 136817 197779 136883 197782
rect 140865 197779 140931 197782
rect 140998 197780 141004 197782
rect 141068 197780 141074 197844
rect 157006 197780 157012 197844
rect 157076 197842 157082 197844
rect 160829 197842 160895 197845
rect 157076 197840 160895 197842
rect 157076 197784 160834 197840
rect 160890 197784 160895 197840
rect 157076 197782 160895 197784
rect 157076 197780 157082 197782
rect 160829 197779 160895 197782
rect 163221 197842 163287 197845
rect 163998 197842 164004 197844
rect 163221 197840 164004 197842
rect 163221 197784 163226 197840
rect 163282 197784 164004 197840
rect 163221 197782 164004 197784
rect 163221 197779 163287 197782
rect 163998 197780 164004 197782
rect 164068 197780 164074 197844
rect 583520 197828 584960 197918
rect 124765 197706 124831 197709
rect 133505 197706 133571 197709
rect 146201 197706 146267 197709
rect 124765 197704 133571 197706
rect 124765 197648 124770 197704
rect 124826 197648 133510 197704
rect 133566 197648 133571 197704
rect 124765 197646 133571 197648
rect 124765 197643 124831 197646
rect 133505 197643 133571 197646
rect 137970 197704 146267 197706
rect 137970 197648 146206 197704
rect 146262 197648 146267 197704
rect 137970 197646 146267 197648
rect 125501 197570 125567 197573
rect 137970 197570 138030 197646
rect 146201 197643 146267 197646
rect 151721 197706 151787 197709
rect 167637 197706 167703 197709
rect 151721 197704 167703 197706
rect 151721 197648 151726 197704
rect 151782 197648 167642 197704
rect 167698 197648 167703 197704
rect 151721 197646 167703 197648
rect 151721 197643 151787 197646
rect 167637 197643 167703 197646
rect 168097 197706 168163 197709
rect 168230 197706 168236 197708
rect 168097 197704 168236 197706
rect 168097 197648 168102 197704
rect 168158 197648 168236 197704
rect 168097 197646 168236 197648
rect 168097 197643 168163 197646
rect 168230 197644 168236 197646
rect 168300 197644 168306 197708
rect 125501 197568 138030 197570
rect 125501 197512 125506 197568
rect 125562 197512 138030 197568
rect 125501 197510 138030 197512
rect 138289 197570 138355 197573
rect 145230 197570 145236 197572
rect 138289 197568 145236 197570
rect 138289 197512 138294 197568
rect 138350 197512 145236 197568
rect 138289 197510 145236 197512
rect 125501 197507 125567 197510
rect 138289 197507 138355 197510
rect 145230 197508 145236 197510
rect 145300 197508 145306 197572
rect 169702 197508 169708 197572
rect 169772 197570 169778 197572
rect 170857 197570 170923 197573
rect 169772 197568 170923 197570
rect 169772 197512 170862 197568
rect 170918 197512 170923 197568
rect 169772 197510 170923 197512
rect 169772 197508 169778 197510
rect 170857 197507 170923 197510
rect 171358 197508 171364 197572
rect 171428 197570 171434 197572
rect 189993 197570 190059 197573
rect 171428 197568 190059 197570
rect 171428 197512 189998 197568
rect 190054 197512 190059 197568
rect 171428 197510 190059 197512
rect 171428 197508 171434 197510
rect 189993 197507 190059 197510
rect 122833 197434 122899 197437
rect 124121 197434 124187 197437
rect 122833 197432 124187 197434
rect -960 197298 480 197388
rect 122833 197376 122838 197432
rect 122894 197376 124126 197432
rect 124182 197376 124187 197432
rect 122833 197374 124187 197376
rect 122833 197371 122899 197374
rect 124121 197371 124187 197374
rect 128997 197434 129063 197437
rect 136817 197434 136883 197437
rect 128997 197432 136883 197434
rect 128997 197376 129002 197432
rect 129058 197376 136822 197432
rect 136878 197376 136883 197432
rect 128997 197374 136883 197376
rect 128997 197371 129063 197374
rect 136817 197371 136883 197374
rect 138933 197434 138999 197437
rect 142470 197434 142476 197436
rect 138933 197432 142476 197434
rect 138933 197376 138938 197432
rect 138994 197376 142476 197432
rect 138933 197374 142476 197376
rect 138933 197371 138999 197374
rect 142470 197372 142476 197374
rect 142540 197372 142546 197436
rect 150525 197434 150591 197437
rect 151118 197434 151124 197436
rect 150525 197432 151124 197434
rect 150525 197376 150530 197432
rect 150586 197376 151124 197432
rect 150525 197374 151124 197376
rect 150525 197371 150591 197374
rect 151118 197372 151124 197374
rect 151188 197372 151194 197436
rect 159265 197434 159331 197437
rect 162025 197434 162091 197437
rect 165889 197434 165955 197437
rect 170765 197436 170831 197437
rect 170765 197434 170812 197436
rect 159265 197432 165955 197434
rect 159265 197376 159270 197432
rect 159326 197376 162030 197432
rect 162086 197376 165894 197432
rect 165950 197376 165955 197432
rect 159265 197374 165955 197376
rect 170720 197432 170812 197434
rect 170720 197376 170770 197432
rect 170720 197374 170812 197376
rect 159265 197371 159331 197374
rect 162025 197371 162091 197374
rect 165889 197371 165955 197374
rect 170765 197372 170812 197374
rect 170876 197372 170882 197436
rect 175733 197434 175799 197437
rect 176510 197434 176516 197436
rect 175733 197432 176516 197434
rect 175733 197376 175738 197432
rect 175794 197376 176516 197432
rect 175733 197374 176516 197376
rect 170765 197371 170831 197372
rect 175733 197371 175799 197374
rect 176510 197372 176516 197374
rect 176580 197372 176586 197436
rect 3141 197298 3207 197301
rect -960 197296 3207 197298
rect -960 197240 3146 197296
rect 3202 197240 3207 197296
rect -960 197238 3207 197240
rect -960 197148 480 197238
rect 3141 197235 3207 197238
rect 131757 197298 131823 197301
rect 132309 197298 132375 197301
rect 580257 197298 580323 197301
rect 131757 197296 580323 197298
rect 131757 197240 131762 197296
rect 131818 197240 132314 197296
rect 132370 197240 580262 197296
rect 580318 197240 580323 197296
rect 131757 197238 580323 197240
rect 131757 197235 131823 197238
rect 132309 197235 132375 197238
rect 580257 197235 580323 197238
rect 125409 197162 125475 197165
rect 131849 197162 131915 197165
rect 125409 197160 131915 197162
rect 125409 197104 125414 197160
rect 125470 197104 131854 197160
rect 131910 197104 131915 197160
rect 125409 197102 131915 197104
rect 125409 197099 125475 197102
rect 131849 197099 131915 197102
rect 132534 197100 132540 197164
rect 132604 197162 132610 197164
rect 133638 197162 133644 197164
rect 132604 197102 133644 197162
rect 132604 197100 132610 197102
rect 133638 197100 133644 197102
rect 133708 197100 133714 197164
rect 140998 197100 141004 197164
rect 141068 197162 141074 197164
rect 141969 197162 142035 197165
rect 141068 197160 142035 197162
rect 141068 197104 141974 197160
rect 142030 197104 142035 197160
rect 141068 197102 142035 197104
rect 141068 197100 141074 197102
rect 141969 197099 142035 197102
rect 144126 197100 144132 197164
rect 144196 197162 144202 197164
rect 144361 197162 144427 197165
rect 144196 197160 144427 197162
rect 144196 197104 144366 197160
rect 144422 197104 144427 197160
rect 144196 197102 144427 197104
rect 144196 197100 144202 197102
rect 144361 197099 144427 197102
rect 146109 197162 146175 197165
rect 147438 197162 147444 197164
rect 146109 197160 147444 197162
rect 146109 197104 146114 197160
rect 146170 197104 147444 197160
rect 146109 197102 147444 197104
rect 146109 197099 146175 197102
rect 147438 197100 147444 197102
rect 147508 197162 147514 197164
rect 445017 197162 445083 197165
rect 147508 197160 445083 197162
rect 147508 197104 445022 197160
rect 445078 197104 445083 197160
rect 147508 197102 445083 197104
rect 147508 197100 147514 197102
rect 445017 197099 445083 197102
rect 62113 197026 62179 197029
rect 159265 197026 159331 197029
rect 62113 197024 159331 197026
rect 62113 196968 62118 197024
rect 62174 196968 159270 197024
rect 159326 196968 159331 197024
rect 62113 196966 159331 196968
rect 62113 196963 62179 196966
rect 159265 196963 159331 196966
rect 163497 197026 163563 197029
rect 173341 197028 173407 197029
rect 163998 197026 164004 197028
rect 163497 197024 164004 197026
rect 163497 196968 163502 197024
rect 163558 196968 164004 197024
rect 163497 196966 164004 196968
rect 163497 196963 163563 196966
rect 163998 196964 164004 196966
rect 164068 196964 164074 197028
rect 173341 197024 173388 197028
rect 173452 197026 173458 197028
rect 177389 197026 177455 197029
rect 210366 197026 210372 197028
rect 173341 196968 173346 197024
rect 173341 196964 173388 196968
rect 173452 196966 173498 197026
rect 177389 197024 210372 197026
rect 177389 196968 177394 197024
rect 177450 196968 210372 197024
rect 177389 196966 210372 196968
rect 173452 196964 173458 196966
rect 173341 196963 173407 196964
rect 177389 196963 177455 196966
rect 210366 196964 210372 196966
rect 210436 197026 210442 197028
rect 210918 197026 210924 197028
rect 210436 196966 210924 197026
rect 210436 196964 210442 196966
rect 210918 196964 210924 196966
rect 210988 196964 210994 197028
rect 105537 196890 105603 196893
rect 170765 196890 170831 196893
rect 420913 196890 420979 196893
rect 105537 196888 170831 196890
rect 105537 196832 105542 196888
rect 105598 196832 170770 196888
rect 170826 196832 170831 196888
rect 105537 196830 170831 196832
rect 105537 196827 105603 196830
rect 170765 196827 170831 196830
rect 209730 196888 420979 196890
rect 209730 196832 420918 196888
rect 420974 196832 420979 196888
rect 209730 196830 420979 196832
rect 122230 196692 122236 196756
rect 122300 196754 122306 196756
rect 135069 196754 135135 196757
rect 122300 196752 135135 196754
rect 122300 196696 135074 196752
rect 135130 196696 135135 196752
rect 122300 196694 135135 196696
rect 122300 196692 122306 196694
rect 135069 196691 135135 196694
rect 138197 196756 138263 196757
rect 138197 196752 138244 196756
rect 138308 196754 138314 196756
rect 138197 196696 138202 196752
rect 138197 196692 138244 196696
rect 138308 196694 138354 196754
rect 138308 196692 138314 196694
rect 139894 196692 139900 196756
rect 139964 196754 139970 196756
rect 140497 196754 140563 196757
rect 139964 196752 140563 196754
rect 139964 196696 140502 196752
rect 140558 196696 140563 196752
rect 139964 196694 140563 196696
rect 139964 196692 139970 196694
rect 138197 196691 138263 196692
rect 140497 196691 140563 196694
rect 143206 196692 143212 196756
rect 143276 196754 143282 196756
rect 143349 196754 143415 196757
rect 149145 196756 149211 196757
rect 149094 196754 149100 196756
rect 143276 196752 143415 196754
rect 143276 196696 143354 196752
rect 143410 196696 143415 196752
rect 143276 196694 143415 196696
rect 149054 196694 149100 196754
rect 149164 196752 149211 196756
rect 149206 196696 149211 196752
rect 143276 196692 143282 196694
rect 143349 196691 143415 196694
rect 149094 196692 149100 196694
rect 149164 196692 149211 196696
rect 149145 196691 149211 196692
rect 151077 196754 151143 196757
rect 151854 196754 151860 196756
rect 151077 196752 151860 196754
rect 151077 196696 151082 196752
rect 151138 196696 151860 196752
rect 151077 196694 151860 196696
rect 151077 196691 151143 196694
rect 151854 196692 151860 196694
rect 151924 196692 151930 196756
rect 156505 196754 156571 196757
rect 161197 196756 161263 196757
rect 157190 196754 157196 196756
rect 156505 196752 157196 196754
rect 156505 196696 156510 196752
rect 156566 196696 157196 196752
rect 156505 196694 157196 196696
rect 156505 196691 156571 196694
rect 157190 196692 157196 196694
rect 157260 196692 157266 196756
rect 161197 196752 161244 196756
rect 161308 196754 161314 196756
rect 163681 196754 163747 196757
rect 163814 196754 163820 196756
rect 161197 196696 161202 196752
rect 161197 196692 161244 196696
rect 161308 196694 161354 196754
rect 163681 196752 163820 196754
rect 163681 196696 163686 196752
rect 163742 196696 163820 196752
rect 163681 196694 163820 196696
rect 161308 196692 161314 196694
rect 161197 196691 161263 196692
rect 163681 196691 163747 196694
rect 163814 196692 163820 196694
rect 163884 196692 163890 196756
rect 164366 196692 164372 196756
rect 164436 196754 164442 196756
rect 164693 196754 164759 196757
rect 164436 196752 164759 196754
rect 164436 196696 164698 196752
rect 164754 196696 164759 196752
rect 164436 196694 164759 196696
rect 164436 196692 164442 196694
rect 164693 196691 164759 196694
rect 170857 196754 170923 196757
rect 170990 196754 170996 196756
rect 170857 196752 170996 196754
rect 170857 196696 170862 196752
rect 170918 196696 170996 196752
rect 170857 196694 170996 196696
rect 170857 196691 170923 196694
rect 170990 196692 170996 196694
rect 171060 196692 171066 196756
rect 173065 196754 173131 196757
rect 205582 196754 205588 196756
rect 173065 196752 205588 196754
rect 173065 196696 173070 196752
rect 173126 196696 205588 196752
rect 173065 196694 205588 196696
rect 173065 196691 173131 196694
rect 205582 196692 205588 196694
rect 205652 196754 205658 196756
rect 209730 196754 209790 196830
rect 420913 196827 420979 196830
rect 205652 196694 209790 196754
rect 205652 196692 205658 196694
rect 210918 196692 210924 196756
rect 210988 196754 210994 196756
rect 576117 196754 576183 196757
rect 210988 196752 576183 196754
rect 210988 196696 576122 196752
rect 576178 196696 576183 196752
rect 210988 196694 576183 196696
rect 210988 196692 210994 196694
rect 576117 196691 576183 196694
rect 117078 196556 117084 196620
rect 117148 196618 117154 196620
rect 146109 196618 146175 196621
rect 117148 196616 146175 196618
rect 117148 196560 146114 196616
rect 146170 196560 146175 196616
rect 117148 196558 146175 196560
rect 117148 196556 117154 196558
rect 146109 196555 146175 196558
rect 146937 196618 147003 196621
rect 149462 196618 149468 196620
rect 146937 196616 149468 196618
rect 146937 196560 146942 196616
rect 146998 196560 149468 196616
rect 146937 196558 149468 196560
rect 146937 196555 147003 196558
rect 149462 196556 149468 196558
rect 149532 196556 149538 196620
rect 164233 196618 164299 196621
rect 190494 196618 190500 196620
rect 164233 196616 190500 196618
rect 164233 196560 164238 196616
rect 164294 196560 190500 196616
rect 164233 196558 190500 196560
rect 164233 196555 164299 196558
rect 190494 196556 190500 196558
rect 190564 196618 190570 196620
rect 576301 196618 576367 196621
rect 190564 196616 576367 196618
rect 190564 196560 576306 196616
rect 576362 196560 576367 196616
rect 190564 196558 576367 196560
rect 190564 196556 190570 196558
rect 576301 196555 576367 196558
rect 132585 196482 132651 196485
rect 133822 196482 133828 196484
rect 132585 196480 133828 196482
rect 132585 196424 132590 196480
rect 132646 196424 133828 196480
rect 132585 196422 133828 196424
rect 132585 196419 132651 196422
rect 133822 196420 133828 196422
rect 133892 196482 133898 196484
rect 137870 196482 137876 196484
rect 133892 196422 137876 196482
rect 133892 196420 133898 196422
rect 137870 196420 137876 196422
rect 137940 196420 137946 196484
rect 138790 196420 138796 196484
rect 138860 196482 138866 196484
rect 141233 196482 141299 196485
rect 138860 196480 141299 196482
rect 138860 196424 141238 196480
rect 141294 196424 141299 196480
rect 138860 196422 141299 196424
rect 138860 196420 138866 196422
rect 141233 196419 141299 196422
rect 148225 196482 148291 196485
rect 153285 196482 153351 196485
rect 148225 196480 153351 196482
rect 148225 196424 148230 196480
rect 148286 196424 153290 196480
rect 153346 196424 153351 196480
rect 148225 196422 153351 196424
rect 148225 196419 148291 196422
rect 153285 196419 153351 196422
rect 156229 196482 156295 196485
rect 157374 196482 157380 196484
rect 156229 196480 157380 196482
rect 156229 196424 156234 196480
rect 156290 196424 157380 196480
rect 156229 196422 157380 196424
rect 156229 196419 156295 196422
rect 157374 196420 157380 196422
rect 157444 196420 157450 196484
rect 169661 196482 169727 196485
rect 171726 196482 171732 196484
rect 169661 196480 171732 196482
rect 169661 196424 169666 196480
rect 169722 196424 171732 196480
rect 169661 196422 171732 196424
rect 169661 196419 169727 196422
rect 171726 196420 171732 196422
rect 171796 196420 171802 196484
rect 172973 196482 173039 196485
rect 198825 196482 198891 196485
rect 172973 196480 198891 196482
rect 172973 196424 172978 196480
rect 173034 196424 198830 196480
rect 198886 196424 198891 196480
rect 172973 196422 198891 196424
rect 172973 196419 173039 196422
rect 198825 196419 198891 196422
rect 132401 196346 132467 196349
rect 135110 196346 135116 196348
rect 132401 196344 135116 196346
rect 132401 196288 132406 196344
rect 132462 196288 135116 196344
rect 132401 196286 135116 196288
rect 132401 196283 132467 196286
rect 135110 196284 135116 196286
rect 135180 196284 135186 196348
rect 167310 196284 167316 196348
rect 167380 196346 167386 196348
rect 168097 196346 168163 196349
rect 167380 196344 168163 196346
rect 167380 196288 168102 196344
rect 168158 196288 168163 196344
rect 167380 196286 168163 196288
rect 167380 196284 167386 196286
rect 168097 196283 168163 196286
rect 137369 196212 137435 196213
rect 137318 196210 137324 196212
rect 137278 196150 137324 196210
rect 137388 196208 137435 196212
rect 137430 196152 137435 196208
rect 137318 196148 137324 196150
rect 137388 196148 137435 196152
rect 137870 196148 137876 196212
rect 137940 196210 137946 196212
rect 138381 196210 138447 196213
rect 137940 196208 138447 196210
rect 137940 196152 138386 196208
rect 138442 196152 138447 196208
rect 137940 196150 138447 196152
rect 137940 196148 137946 196150
rect 137369 196147 137435 196148
rect 138381 196147 138447 196150
rect 153285 196210 153351 196213
rect 154062 196210 154068 196212
rect 153285 196208 154068 196210
rect 153285 196152 153290 196208
rect 153346 196152 154068 196208
rect 153285 196150 154068 196152
rect 153285 196147 153351 196150
rect 154062 196148 154068 196150
rect 154132 196148 154138 196212
rect 136633 196074 136699 196077
rect 152641 196076 152707 196077
rect 139342 196074 139348 196076
rect 136633 196072 139348 196074
rect 136633 196016 136638 196072
rect 136694 196016 139348 196072
rect 136633 196014 139348 196016
rect 136633 196011 136699 196014
rect 139342 196012 139348 196014
rect 139412 196012 139418 196076
rect 152590 196012 152596 196076
rect 152660 196074 152707 196076
rect 153377 196074 153443 196077
rect 153878 196074 153884 196076
rect 152660 196072 152752 196074
rect 152702 196016 152752 196072
rect 152660 196014 152752 196016
rect 153377 196072 153884 196074
rect 153377 196016 153382 196072
rect 153438 196016 153884 196072
rect 153377 196014 153884 196016
rect 152660 196012 152707 196014
rect 152641 196011 152707 196012
rect 153377 196011 153443 196014
rect 153878 196012 153884 196014
rect 153948 196012 153954 196076
rect 154246 196012 154252 196076
rect 154316 196074 154322 196076
rect 154481 196074 154547 196077
rect 154316 196072 154547 196074
rect 154316 196016 154486 196072
rect 154542 196016 154547 196072
rect 154316 196014 154547 196016
rect 154316 196012 154322 196014
rect 154481 196011 154547 196014
rect 156413 196074 156479 196077
rect 156638 196074 156644 196076
rect 156413 196072 156644 196074
rect 156413 196016 156418 196072
rect 156474 196016 156644 196072
rect 156413 196014 156644 196016
rect 156413 196011 156479 196014
rect 156638 196012 156644 196014
rect 156708 196012 156714 196076
rect 174537 196074 174603 196077
rect 174670 196074 174676 196076
rect 174537 196072 174676 196074
rect 174537 196016 174542 196072
rect 174598 196016 174676 196072
rect 174537 196014 174676 196016
rect 174537 196011 174603 196014
rect 174670 196012 174676 196014
rect 174740 196012 174746 196076
rect 122598 195876 122604 195940
rect 122668 195938 122674 195940
rect 122833 195938 122899 195941
rect 122668 195936 122899 195938
rect 122668 195880 122838 195936
rect 122894 195880 122899 195936
rect 122668 195878 122899 195880
rect 122668 195876 122674 195878
rect 122833 195875 122899 195878
rect 136030 195876 136036 195940
rect 136100 195938 136106 195940
rect 136173 195938 136239 195941
rect 136449 195940 136515 195941
rect 136100 195936 136239 195938
rect 136100 195880 136178 195936
rect 136234 195880 136239 195936
rect 136100 195878 136239 195880
rect 136100 195876 136106 195878
rect 136173 195875 136239 195878
rect 136398 195876 136404 195940
rect 136468 195938 136515 195940
rect 136725 195938 136791 195941
rect 138381 195940 138447 195941
rect 137134 195938 137140 195940
rect 136468 195936 136560 195938
rect 136510 195880 136560 195936
rect 136468 195878 136560 195880
rect 136725 195936 137140 195938
rect 136725 195880 136730 195936
rect 136786 195880 137140 195936
rect 136725 195878 137140 195880
rect 136468 195876 136515 195878
rect 136449 195875 136515 195876
rect 136725 195875 136791 195878
rect 137134 195876 137140 195878
rect 137204 195876 137210 195940
rect 138381 195938 138428 195940
rect 138336 195936 138428 195938
rect 138336 195880 138386 195936
rect 138336 195878 138428 195880
rect 138381 195876 138428 195878
rect 138492 195876 138498 195940
rect 138606 195876 138612 195940
rect 138676 195938 138682 195940
rect 139117 195938 139183 195941
rect 138676 195936 139183 195938
rect 138676 195880 139122 195936
rect 139178 195880 139183 195936
rect 138676 195878 139183 195880
rect 138676 195876 138682 195878
rect 138381 195875 138447 195876
rect 139117 195875 139183 195878
rect 143165 195938 143231 195941
rect 143942 195938 143948 195940
rect 143165 195936 143948 195938
rect 143165 195880 143170 195936
rect 143226 195880 143948 195936
rect 143165 195878 143948 195880
rect 143165 195875 143231 195878
rect 143942 195876 143948 195878
rect 144012 195938 144018 195940
rect 485773 195938 485839 195941
rect 144012 195936 485839 195938
rect 144012 195880 485778 195936
rect 485834 195880 485839 195936
rect 144012 195878 485839 195880
rect 144012 195876 144018 195878
rect 485773 195875 485839 195878
rect 102961 195802 103027 195805
rect 173433 195802 173499 195805
rect 102961 195800 173499 195802
rect 102961 195744 102966 195800
rect 103022 195744 173438 195800
rect 173494 195744 173499 195800
rect 102961 195742 173499 195744
rect 102961 195739 103027 195742
rect 173433 195739 173499 195742
rect 174721 195802 174787 195805
rect 174854 195802 174860 195804
rect 174721 195800 174860 195802
rect 174721 195744 174726 195800
rect 174782 195744 174860 195800
rect 174721 195742 174860 195744
rect 174721 195739 174787 195742
rect 174854 195740 174860 195742
rect 174924 195740 174930 195804
rect 212441 195802 212507 195805
rect 386413 195802 386479 195805
rect 212441 195800 386479 195802
rect 212441 195744 212446 195800
rect 212502 195744 386418 195800
rect 386474 195744 386479 195800
rect 212441 195742 386479 195744
rect 212441 195739 212507 195742
rect 386413 195739 386479 195742
rect 124070 195604 124076 195668
rect 124140 195666 124146 195668
rect 134885 195666 134951 195669
rect 124140 195664 134951 195666
rect 124140 195608 134890 195664
rect 134946 195608 134951 195664
rect 124140 195606 134951 195608
rect 124140 195604 124146 195606
rect 134885 195603 134951 195606
rect 170949 195666 171015 195669
rect 211521 195666 211587 195669
rect 220077 195666 220143 195669
rect 170949 195664 220143 195666
rect 170949 195608 170954 195664
rect 171010 195608 211526 195664
rect 211582 195608 220082 195664
rect 220138 195608 220143 195664
rect 170949 195606 220143 195608
rect 170949 195603 171015 195606
rect 211521 195603 211587 195606
rect 220077 195603 220143 195606
rect 130561 195530 130627 195533
rect 143993 195530 144059 195533
rect 130561 195528 144059 195530
rect 130561 195472 130566 195528
rect 130622 195472 143998 195528
rect 144054 195472 144059 195528
rect 130561 195470 144059 195472
rect 130561 195467 130627 195470
rect 143993 195467 144059 195470
rect 153837 195530 153903 195533
rect 218053 195530 218119 195533
rect 582833 195530 582899 195533
rect 153837 195528 582899 195530
rect 153837 195472 153842 195528
rect 153898 195472 218058 195528
rect 218114 195472 582838 195528
rect 582894 195472 582899 195528
rect 153837 195470 582899 195472
rect 153837 195467 153903 195470
rect 218053 195467 218119 195470
rect 582833 195467 582899 195470
rect 104709 195394 104775 195397
rect 136633 195394 136699 195397
rect 164509 195396 164575 195397
rect 164509 195394 164556 195396
rect 104709 195392 136699 195394
rect 104709 195336 104714 195392
rect 104770 195336 136638 195392
rect 136694 195336 136699 195392
rect 104709 195334 136699 195336
rect 164464 195392 164556 195394
rect 164464 195336 164514 195392
rect 164464 195334 164556 195336
rect 104709 195331 104775 195334
rect 136633 195331 136699 195334
rect 164509 195332 164556 195334
rect 164620 195332 164626 195396
rect 165470 195332 165476 195396
rect 165540 195394 165546 195396
rect 194593 195394 194659 195397
rect 571977 195394 572043 195397
rect 165540 195392 572043 195394
rect 165540 195336 194598 195392
rect 194654 195336 571982 195392
rect 572038 195336 572043 195392
rect 165540 195334 572043 195336
rect 165540 195332 165546 195334
rect 164509 195331 164575 195332
rect 194593 195331 194659 195334
rect 571977 195331 572043 195334
rect 96337 195258 96403 195261
rect 165429 195258 165495 195261
rect 168598 195258 168604 195260
rect 96337 195256 168604 195258
rect 96337 195200 96342 195256
rect 96398 195200 165434 195256
rect 165490 195200 168604 195256
rect 96337 195198 168604 195200
rect 96337 195195 96403 195198
rect 165429 195195 165495 195198
rect 168598 195196 168604 195198
rect 168668 195196 168674 195260
rect 189073 195258 189139 195261
rect 189901 195258 189967 195261
rect 577497 195258 577563 195261
rect 189073 195256 577563 195258
rect 189073 195200 189078 195256
rect 189134 195200 189906 195256
rect 189962 195200 577502 195256
rect 577558 195200 577563 195256
rect 189073 195198 577563 195200
rect 189073 195195 189139 195198
rect 189901 195195 189967 195198
rect 577497 195195 577563 195198
rect 142981 195124 143047 195125
rect 142981 195122 143028 195124
rect 142936 195120 143028 195122
rect 142936 195064 142986 195120
rect 142936 195062 143028 195064
rect 142981 195060 143028 195062
rect 143092 195060 143098 195124
rect 181805 195122 181871 195125
rect 214046 195122 214052 195124
rect 181805 195120 214052 195122
rect 181805 195064 181810 195120
rect 181866 195064 214052 195120
rect 181805 195062 214052 195064
rect 142981 195059 143047 195060
rect 181805 195059 181871 195062
rect 214046 195060 214052 195062
rect 214116 195122 214122 195124
rect 558913 195122 558979 195125
rect 214116 195120 558979 195122
rect 214116 195064 558918 195120
rect 558974 195064 558979 195120
rect 214116 195062 558979 195064
rect 214116 195060 214122 195062
rect 558913 195059 558979 195062
rect 170213 194986 170279 194989
rect 211153 194986 211219 194989
rect 212441 194986 212507 194989
rect 170213 194984 212507 194986
rect 170213 194928 170218 194984
rect 170274 194928 211158 194984
rect 211214 194928 212446 194984
rect 212502 194928 212507 194984
rect 170213 194926 212507 194928
rect 170213 194923 170279 194926
rect 211153 194923 211219 194926
rect 212441 194923 212507 194926
rect 171409 194850 171475 194853
rect 189073 194850 189139 194853
rect 171409 194848 189139 194850
rect 171409 194792 171414 194848
rect 171470 194792 189078 194848
rect 189134 194792 189139 194848
rect 171409 194790 189139 194792
rect 171409 194787 171475 194790
rect 189073 194787 189139 194790
rect 121361 194580 121427 194581
rect 121310 194578 121316 194580
rect 121270 194518 121316 194578
rect 121380 194576 121427 194580
rect 121422 194520 121427 194576
rect 121310 194516 121316 194518
rect 121380 194516 121427 194520
rect 121361 194515 121427 194516
rect 144177 194578 144243 194581
rect 145005 194578 145071 194581
rect 144177 194576 145071 194578
rect 144177 194520 144182 194576
rect 144238 194520 145010 194576
rect 145066 194520 145071 194576
rect 144177 194518 145071 194520
rect 144177 194515 144243 194518
rect 145005 194515 145071 194518
rect 152641 194578 152707 194581
rect 542353 194578 542419 194581
rect 152641 194576 542419 194578
rect 152641 194520 152646 194576
rect 152702 194520 542358 194576
rect 542414 194520 542419 194576
rect 152641 194518 542419 194520
rect 152641 194515 152707 194518
rect 542353 194515 542419 194518
rect 425053 194442 425119 194445
rect 144870 194440 425119 194442
rect 144870 194384 425058 194440
rect 425114 194384 425119 194440
rect 144870 194382 425119 194384
rect 126973 194306 127039 194309
rect 134701 194306 134767 194309
rect 126973 194304 134767 194306
rect 126973 194248 126978 194304
rect 127034 194248 134706 194304
rect 134762 194248 134767 194304
rect 126973 194246 134767 194248
rect 126973 194243 127039 194246
rect 134701 194243 134767 194246
rect 108798 194108 108804 194172
rect 108868 194170 108874 194172
rect 142286 194170 142292 194172
rect 108868 194110 142292 194170
rect 108868 194108 108874 194110
rect 142286 194108 142292 194110
rect 142356 194170 142362 194172
rect 144870 194170 144930 194382
rect 425053 194379 425119 194382
rect 147121 194306 147187 194309
rect 340873 194306 340939 194309
rect 147121 194304 340939 194306
rect 147121 194248 147126 194304
rect 147182 194248 340878 194304
rect 340934 194248 340939 194304
rect 147121 194246 340939 194248
rect 147121 194243 147187 194246
rect 340873 194243 340939 194246
rect 142356 194110 144930 194170
rect 178585 194170 178651 194173
rect 202229 194170 202295 194173
rect 178585 194168 202295 194170
rect 178585 194112 178590 194168
rect 178646 194112 202234 194168
rect 202290 194112 202295 194168
rect 178585 194110 202295 194112
rect 142356 194108 142362 194110
rect 178585 194107 178651 194110
rect 202229 194107 202295 194110
rect 88977 194034 89043 194037
rect 99230 194034 99236 194036
rect 88977 194032 99236 194034
rect 88977 193976 88982 194032
rect 89038 193976 99236 194032
rect 88977 193974 99236 193976
rect 88977 193971 89043 193974
rect 99230 193972 99236 193974
rect 99300 194034 99306 194036
rect 152273 194034 152339 194037
rect 99300 194032 152339 194034
rect 99300 193976 152278 194032
rect 152334 193976 152339 194032
rect 99300 193974 152339 193976
rect 99300 193972 99306 193974
rect 152273 193971 152339 193974
rect 197302 193972 197308 194036
rect 197372 194034 197378 194036
rect 237373 194034 237439 194037
rect 581729 194034 581795 194037
rect 197372 194032 237439 194034
rect 197372 193976 237378 194032
rect 237434 193976 237439 194032
rect 197372 193974 237439 193976
rect 197372 193972 197378 193974
rect 237373 193971 237439 193974
rect 567150 194032 581795 194034
rect 567150 193976 581734 194032
rect 581790 193976 581795 194032
rect 567150 193974 581795 193976
rect 27613 193898 27679 193901
rect 119654 193898 119660 193900
rect 27613 193896 119660 193898
rect 27613 193840 27618 193896
rect 27674 193840 119660 193896
rect 27613 193838 119660 193840
rect 27613 193835 27679 193838
rect 119654 193836 119660 193838
rect 119724 193836 119730 193900
rect 123477 193898 123543 193901
rect 128905 193898 128971 193901
rect 123477 193896 128971 193898
rect 123477 193840 123482 193896
rect 123538 193840 128910 193896
rect 128966 193840 128971 193896
rect 123477 193838 128971 193840
rect 123477 193835 123543 193838
rect 128905 193835 128971 193838
rect 168005 193898 168071 193901
rect 198774 193898 198780 193900
rect 168005 193896 198780 193898
rect 168005 193840 168010 193896
rect 168066 193840 198780 193896
rect 168005 193838 198780 193840
rect 168005 193835 168071 193838
rect 198774 193836 198780 193838
rect 198844 193898 198850 193900
rect 567150 193898 567210 193974
rect 581729 193971 581795 193974
rect 198844 193838 567210 193898
rect 579797 193898 579863 193901
rect 583520 193898 584960 193988
rect 579797 193896 584960 193898
rect 579797 193840 579802 193896
rect 579858 193840 584960 193896
rect 579797 193838 584960 193840
rect 198844 193836 198850 193838
rect 579797 193835 579863 193838
rect 146661 193764 146727 193765
rect 154113 193764 154179 193765
rect 146661 193762 146708 193764
rect 146616 193760 146708 193762
rect 146616 193704 146666 193760
rect 146616 193702 146708 193704
rect 146661 193700 146708 193702
rect 146772 193700 146778 193764
rect 154062 193762 154068 193764
rect 154022 193702 154068 193762
rect 154132 193760 154179 193764
rect 154174 193704 154179 193760
rect 583520 193748 584960 193838
rect 154062 193700 154068 193702
rect 154132 193700 154179 193704
rect 146661 193699 146727 193700
rect 154113 193699 154179 193700
rect -960 193218 480 193308
rect 134190 193292 134196 193356
rect 134260 193354 134266 193356
rect 134333 193354 134399 193357
rect 134260 193352 134399 193354
rect 134260 193296 134338 193352
rect 134394 193296 134399 193352
rect 134260 193294 134399 193296
rect 134260 193292 134266 193294
rect 134333 193291 134399 193294
rect 3417 193218 3483 193221
rect -960 193216 3483 193218
rect -960 193160 3422 193216
rect 3478 193160 3483 193216
rect -960 193158 3483 193160
rect -960 193068 480 193158
rect 3417 193155 3483 193158
rect 34513 193218 34579 193221
rect 172513 193218 172579 193221
rect 173709 193218 173775 193221
rect 34513 193216 173775 193218
rect 34513 193160 34518 193216
rect 34574 193160 172518 193216
rect 172574 193160 173714 193216
rect 173770 193160 173775 193216
rect 34513 193158 173775 193160
rect 34513 193155 34579 193158
rect 172513 193155 172579 193158
rect 173709 193155 173775 193158
rect 175222 193156 175228 193220
rect 175292 193218 175298 193220
rect 176377 193218 176443 193221
rect 175292 193216 176443 193218
rect 175292 193160 176382 193216
rect 176438 193160 176443 193216
rect 175292 193158 176443 193160
rect 175292 193156 175298 193158
rect 176377 193155 176443 193158
rect 98637 193082 98703 193085
rect 173014 193082 173020 193084
rect 98637 193080 173020 193082
rect 98637 193024 98642 193080
rect 98698 193024 173020 193080
rect 98637 193022 173020 193024
rect 98637 193019 98703 193022
rect 173014 193020 173020 193022
rect 173084 193082 173090 193084
rect 205766 193082 205772 193084
rect 173084 193022 205772 193082
rect 173084 193020 173090 193022
rect 205766 193020 205772 193022
rect 205836 193020 205842 193084
rect 119654 192884 119660 192948
rect 119724 192946 119730 192948
rect 147581 192946 147647 192949
rect 149094 192946 149100 192948
rect 119724 192886 142170 192946
rect 119724 192884 119730 192886
rect 142110 192810 142170 192886
rect 147581 192944 149100 192946
rect 147581 192888 147586 192944
rect 147642 192888 149100 192944
rect 147581 192886 149100 192888
rect 147581 192883 147647 192886
rect 149094 192884 149100 192886
rect 149164 192884 149170 192948
rect 164366 192884 164372 192948
rect 164436 192946 164442 192948
rect 198825 192946 198891 192949
rect 164436 192944 198891 192946
rect 164436 192888 198830 192944
rect 198886 192888 198891 192944
rect 164436 192886 198891 192888
rect 164436 192884 164442 192886
rect 198825 192883 198891 192886
rect 147489 192810 147555 192813
rect 142110 192808 147555 192810
rect 142110 192752 147494 192808
rect 147550 192752 147555 192808
rect 142110 192750 147555 192752
rect 147489 192747 147555 192750
rect 168414 192748 168420 192812
rect 168484 192810 168490 192812
rect 201585 192810 201651 192813
rect 224217 192810 224283 192813
rect 168484 192808 224283 192810
rect 168484 192752 201590 192808
rect 201646 192752 224222 192808
rect 224278 192752 224283 192808
rect 168484 192750 224283 192752
rect 168484 192748 168490 192750
rect 201585 192747 201651 192750
rect 224217 192747 224283 192750
rect 174721 192674 174787 192677
rect 214097 192674 214163 192677
rect 574829 192674 574895 192677
rect 174721 192672 574895 192674
rect 174721 192616 174726 192672
rect 174782 192616 214102 192672
rect 214158 192616 574834 192672
rect 574890 192616 574895 192672
rect 174721 192614 574895 192616
rect 174721 192611 174787 192614
rect 214097 192611 214163 192614
rect 574829 192611 574895 192614
rect 124029 192538 124095 192541
rect 127893 192538 127959 192541
rect 124029 192536 127959 192538
rect 124029 192480 124034 192536
rect 124090 192480 127898 192536
rect 127954 192480 127959 192536
rect 124029 192478 127959 192480
rect 124029 192475 124095 192478
rect 127893 192475 127959 192478
rect 166390 192476 166396 192540
rect 166460 192538 166466 192540
rect 200614 192538 200620 192540
rect 166460 192478 200620 192538
rect 166460 192476 166466 192478
rect 200614 192476 200620 192478
rect 200684 192538 200690 192540
rect 578233 192538 578299 192541
rect 200684 192536 578299 192538
rect 200684 192480 578238 192536
rect 578294 192480 578299 192536
rect 200684 192478 578299 192480
rect 200684 192476 200690 192478
rect 578233 192475 578299 192478
rect 106917 191722 106983 191725
rect 153142 191722 153148 191724
rect 106917 191720 153148 191722
rect 106917 191664 106922 191720
rect 106978 191664 153148 191720
rect 106917 191662 153148 191664
rect 106917 191659 106983 191662
rect 153142 191660 153148 191662
rect 153212 191722 153218 191724
rect 168833 191722 168899 191725
rect 153212 191720 168899 191722
rect 153212 191664 168838 191720
rect 168894 191664 168899 191720
rect 153212 191662 168899 191664
rect 153212 191660 153218 191662
rect 168833 191659 168899 191662
rect 150433 191586 150499 191589
rect 113130 191584 150499 191586
rect 113130 191528 150438 191584
rect 150494 191528 150499 191584
rect 113130 191526 150499 191528
rect 97625 191178 97691 191181
rect 111885 191178 111951 191181
rect 113130 191178 113190 191526
rect 150433 191523 150499 191526
rect 167862 191524 167868 191588
rect 167932 191586 167938 191588
rect 202086 191586 202092 191588
rect 167932 191526 202092 191586
rect 167932 191524 167938 191526
rect 202086 191524 202092 191526
rect 202156 191586 202162 191588
rect 416773 191586 416839 191589
rect 202156 191584 416839 191586
rect 202156 191528 416778 191584
rect 416834 191528 416839 191584
rect 202156 191526 416839 191528
rect 202156 191524 202162 191526
rect 416773 191523 416839 191526
rect 182081 191450 182147 191453
rect 440233 191450 440299 191453
rect 182081 191448 440299 191450
rect 182081 191392 182086 191448
rect 182142 191392 440238 191448
rect 440294 191392 440299 191448
rect 182081 191390 440299 191392
rect 182081 191387 182147 191390
rect 440233 191387 440299 191390
rect 166574 191252 166580 191316
rect 166644 191314 166650 191316
rect 201033 191314 201099 191317
rect 516133 191314 516199 191317
rect 166644 191312 516199 191314
rect 166644 191256 201038 191312
rect 201094 191256 516138 191312
rect 516194 191256 516199 191312
rect 166644 191254 516199 191256
rect 166644 191252 166650 191254
rect 201033 191251 201099 191254
rect 516133 191251 516199 191254
rect 97625 191176 113190 191178
rect 97625 191120 97630 191176
rect 97686 191120 111890 191176
rect 111946 191120 113190 191176
rect 97625 191118 113190 191120
rect 119705 191178 119771 191181
rect 122598 191178 122604 191180
rect 119705 191176 122604 191178
rect 119705 191120 119710 191176
rect 119766 191120 122604 191176
rect 119705 191118 122604 191120
rect 97625 191115 97691 191118
rect 111885 191115 111951 191118
rect 119705 191115 119771 191118
rect 122598 191116 122604 191118
rect 122668 191178 122674 191180
rect 155861 191178 155927 191181
rect 122668 191176 155927 191178
rect 122668 191120 155866 191176
rect 155922 191120 155927 191176
rect 122668 191118 155927 191120
rect 122668 191116 122674 191118
rect 155861 191115 155927 191118
rect 156822 191116 156828 191180
rect 156892 191178 156898 191180
rect 182081 191178 182147 191181
rect 156892 191176 182147 191178
rect 156892 191120 182086 191176
rect 182142 191120 182147 191176
rect 156892 191118 182147 191120
rect 156892 191116 156898 191118
rect 182081 191115 182147 191118
rect 187141 191178 187207 191181
rect 567837 191178 567903 191181
rect 187141 191176 567903 191178
rect 187141 191120 187146 191176
rect 187202 191120 567842 191176
rect 567898 191120 567903 191176
rect 187141 191118 567903 191120
rect 187141 191115 187207 191118
rect 567837 191115 567903 191118
rect 89069 191042 89135 191045
rect 114134 191042 114140 191044
rect 89069 191040 114140 191042
rect 89069 190984 89074 191040
rect 89130 190984 114140 191040
rect 89069 190982 114140 190984
rect 89069 190979 89135 190982
rect 114134 190980 114140 190982
rect 114204 191042 114210 191044
rect 148133 191042 148199 191045
rect 114204 191040 148199 191042
rect 114204 190984 148138 191040
rect 148194 190984 148199 191040
rect 114204 190982 148199 190984
rect 114204 190980 114210 190982
rect 148133 190979 148199 190982
rect 161238 190980 161244 191044
rect 161308 191042 161314 191044
rect 179321 191042 179387 191045
rect 576209 191042 576275 191045
rect 161308 191040 576275 191042
rect 161308 190984 179326 191040
rect 179382 190984 576214 191040
rect 576270 190984 576275 191040
rect 161308 190982 576275 190984
rect 161308 190980 161314 190982
rect 179321 190979 179387 190982
rect 576209 190979 576275 190982
rect 166022 190844 166028 190908
rect 166092 190906 166098 190908
rect 187141 190906 187207 190909
rect 166092 190904 187207 190906
rect 166092 190848 187146 190904
rect 187202 190848 187207 190904
rect 166092 190846 187207 190848
rect 166092 190844 166098 190846
rect 187141 190843 187207 190846
rect 173709 190770 173775 190773
rect 189022 190770 189028 190772
rect 173709 190768 189028 190770
rect 173709 190712 173714 190768
rect 173770 190712 189028 190768
rect 173709 190710 189028 190712
rect 173709 190707 173775 190710
rect 189022 190708 189028 190710
rect 189092 190708 189098 190772
rect 163814 190572 163820 190636
rect 163884 190634 163890 190636
rect 197302 190634 197308 190636
rect 163884 190574 197308 190634
rect 163884 190572 163890 190574
rect 197302 190572 197308 190574
rect 197372 190572 197378 190636
rect 113030 190436 113036 190500
rect 113100 190498 113106 190500
rect 133229 190498 133295 190501
rect 113100 190496 133295 190498
rect 113100 190440 133234 190496
rect 133290 190440 133295 190496
rect 113100 190438 133295 190440
rect 113100 190436 113106 190438
rect 133229 190435 133295 190438
rect 137277 190364 137343 190365
rect 137277 190360 137324 190364
rect 137388 190362 137394 190364
rect 137277 190304 137282 190360
rect 137277 190300 137324 190304
rect 137388 190302 137434 190362
rect 137388 190300 137394 190302
rect 148174 190300 148180 190364
rect 148244 190362 148250 190364
rect 574921 190362 574987 190365
rect 148244 190360 574987 190362
rect 148244 190304 574926 190360
rect 574982 190304 574987 190360
rect 148244 190302 574987 190304
rect 148244 190300 148250 190302
rect 137277 190299 137343 190300
rect 574921 190299 574987 190302
rect 12433 190226 12499 190229
rect 175406 190226 175412 190228
rect 12433 190224 175412 190226
rect 12433 190168 12438 190224
rect 12494 190168 175412 190224
rect 12433 190166 175412 190168
rect 12433 190163 12499 190166
rect 175406 190164 175412 190166
rect 175476 190164 175482 190228
rect 163446 190028 163452 190092
rect 163516 190090 163522 190092
rect 191966 190090 191972 190092
rect 163516 190030 191972 190090
rect 163516 190028 163522 190030
rect 191966 190028 191972 190030
rect 192036 190090 192042 190092
rect 193070 190090 193076 190092
rect 192036 190030 193076 190090
rect 192036 190028 192042 190030
rect 193070 190028 193076 190030
rect 193140 190028 193146 190092
rect 187734 189892 187740 189956
rect 187804 189954 187810 189956
rect 371233 189954 371299 189957
rect 187804 189952 371299 189954
rect 187804 189896 371238 189952
rect 371294 189896 371299 189952
rect 187804 189894 371299 189896
rect 187804 189892 187810 189894
rect 371233 189891 371299 189894
rect 119654 189756 119660 189820
rect 119724 189818 119730 189820
rect 152641 189818 152707 189821
rect 119724 189816 152707 189818
rect 119724 189760 152646 189816
rect 152702 189760 152707 189816
rect 119724 189758 152707 189760
rect 119724 189756 119730 189758
rect 152641 189755 152707 189758
rect 172278 189756 172284 189820
rect 172348 189818 172354 189820
rect 214373 189818 214439 189821
rect 566549 189818 566615 189821
rect 172348 189816 566615 189818
rect 172348 189760 214378 189816
rect 214434 189760 566554 189816
rect 566610 189760 566615 189816
rect 172348 189758 566615 189760
rect 172348 189756 172354 189758
rect 214373 189755 214439 189758
rect 566549 189755 566615 189758
rect 579613 189818 579679 189821
rect 583520 189818 584960 189908
rect 579613 189816 584960 189818
rect 579613 189760 579618 189816
rect 579674 189760 584960 189816
rect 579613 189758 584960 189760
rect 579613 189755 579679 189758
rect 118366 189620 118372 189684
rect 118436 189682 118442 189684
rect 152457 189682 152523 189685
rect 118436 189680 152523 189682
rect 118436 189624 152462 189680
rect 152518 189624 152523 189680
rect 118436 189622 152523 189624
rect 118436 189620 118442 189622
rect 152457 189619 152523 189622
rect 153653 189682 153719 189685
rect 187734 189682 187740 189684
rect 153653 189680 187740 189682
rect 153653 189624 153658 189680
rect 153714 189624 187740 189680
rect 153653 189622 187740 189624
rect 153653 189619 153719 189622
rect 187734 189620 187740 189622
rect 187804 189620 187810 189684
rect 193070 189620 193076 189684
rect 193140 189682 193146 189684
rect 575105 189682 575171 189685
rect 193140 189680 575171 189682
rect 193140 189624 575110 189680
rect 575166 189624 575171 189680
rect 583520 189668 584960 189758
rect 193140 189622 575171 189624
rect 193140 189620 193146 189622
rect 575105 189619 575171 189622
rect -960 189138 480 189228
rect 3417 189138 3483 189141
rect -960 189136 3483 189138
rect -960 189080 3422 189136
rect 3478 189080 3483 189136
rect -960 189078 3483 189080
rect -960 188988 480 189078
rect 3417 189075 3483 189078
rect 147305 189138 147371 189141
rect 148174 189138 148180 189140
rect 147305 189136 148180 189138
rect 147305 189080 147310 189136
rect 147366 189080 148180 189136
rect 147305 189078 148180 189080
rect 147305 189075 147371 189078
rect 148174 189076 148180 189078
rect 148244 189076 148250 189140
rect 150893 189138 150959 189141
rect 163589 189140 163655 189141
rect 175457 189140 175523 189141
rect 151118 189138 151124 189140
rect 150893 189136 151124 189138
rect 150893 189080 150898 189136
rect 150954 189080 151124 189136
rect 150893 189078 151124 189080
rect 150893 189075 150959 189078
rect 151118 189076 151124 189078
rect 151188 189076 151194 189140
rect 163589 189136 163636 189140
rect 163700 189138 163706 189140
rect 175406 189138 175412 189140
rect 163589 189080 163594 189136
rect 163589 189076 163636 189080
rect 163700 189078 163746 189138
rect 175366 189078 175412 189138
rect 175476 189136 175523 189140
rect 175518 189080 175523 189136
rect 163700 189076 163706 189078
rect 175406 189076 175412 189078
rect 175476 189076 175523 189080
rect 163589 189075 163655 189076
rect 175457 189075 175523 189076
rect 144494 188940 144500 189004
rect 144564 189002 144570 189004
rect 144637 189002 144703 189005
rect 144564 189000 144703 189002
rect 144564 188944 144642 189000
rect 144698 188944 144703 189000
rect 144564 188942 144703 188944
rect 144564 188940 144570 188942
rect 144637 188939 144703 188942
rect 153561 189002 153627 189005
rect 242157 189002 242223 189005
rect 153561 189000 242223 189002
rect 153561 188944 153566 189000
rect 153622 188944 242162 189000
rect 242218 188944 242223 189000
rect 153561 188942 242223 188944
rect 153561 188939 153627 188942
rect 242157 188939 242223 188942
rect 94497 188866 94563 188869
rect 94497 188864 161490 188866
rect 94497 188808 94502 188864
rect 94558 188808 161490 188864
rect 94497 188806 161490 188808
rect 94497 188803 94563 188806
rect 143441 188732 143507 188733
rect 143390 188730 143396 188732
rect 143350 188670 143396 188730
rect 143460 188728 143507 188732
rect 143502 188672 143507 188728
rect 143390 188668 143396 188670
rect 143460 188668 143507 188672
rect 143441 188667 143507 188668
rect 98821 188594 98887 188597
rect 109033 188594 109099 188597
rect 98821 188592 109099 188594
rect 98821 188536 98826 188592
rect 98882 188536 109038 188592
rect 109094 188536 109099 188592
rect 98821 188534 109099 188536
rect 98821 188531 98887 188534
rect 109033 188531 109099 188534
rect 122414 188532 122420 188596
rect 122484 188594 122490 188596
rect 153561 188594 153627 188597
rect 122484 188592 153627 188594
rect 122484 188536 153566 188592
rect 153622 188536 153627 188592
rect 122484 188534 153627 188536
rect 122484 188532 122490 188534
rect 153561 188531 153627 188534
rect 132534 188458 132540 188460
rect 103470 188398 132540 188458
rect 77937 188322 78003 188325
rect 99189 188322 99255 188325
rect 103470 188322 103530 188398
rect 132534 188396 132540 188398
rect 132604 188396 132610 188460
rect 161430 188458 161490 188806
rect 176510 188532 176516 188596
rect 176580 188594 176586 188596
rect 209037 188594 209103 188597
rect 176580 188592 209790 188594
rect 176580 188536 209042 188592
rect 209098 188536 209790 188592
rect 176580 188534 209790 188536
rect 176580 188532 176586 188534
rect 209037 188531 209103 188534
rect 162526 188458 162532 188460
rect 161430 188398 162532 188458
rect 162526 188396 162532 188398
rect 162596 188458 162602 188460
rect 201534 188458 201540 188460
rect 162596 188398 201540 188458
rect 162596 188396 162602 188398
rect 201534 188396 201540 188398
rect 201604 188396 201610 188460
rect 209730 188458 209790 188534
rect 378133 188458 378199 188461
rect 209730 188456 378199 188458
rect 209730 188400 378138 188456
rect 378194 188400 378199 188456
rect 209730 188398 378199 188400
rect 378133 188395 378199 188398
rect 77937 188320 103530 188322
rect 77937 188264 77942 188320
rect 77998 188264 99194 188320
rect 99250 188264 103530 188320
rect 77937 188262 103530 188264
rect 109033 188322 109099 188325
rect 110137 188322 110203 188325
rect 143574 188322 143580 188324
rect 109033 188320 143580 188322
rect 109033 188264 109038 188320
rect 109094 188264 110142 188320
rect 110198 188264 143580 188320
rect 109033 188262 143580 188264
rect 77937 188259 78003 188262
rect 99189 188259 99255 188262
rect 109033 188259 109099 188262
rect 110137 188259 110203 188262
rect 143574 188260 143580 188262
rect 143644 188260 143650 188324
rect 151486 188260 151492 188324
rect 151556 188322 151562 188324
rect 218513 188322 218579 188325
rect 546493 188322 546559 188325
rect 151556 188320 546559 188322
rect 151556 188264 218518 188320
rect 218574 188264 546498 188320
rect 546554 188264 546559 188320
rect 151556 188262 546559 188264
rect 151556 188260 151562 188262
rect 218513 188259 218579 188262
rect 546493 188259 546559 188262
rect 42793 187642 42859 187645
rect 169702 187642 169708 187644
rect 42793 187640 169708 187642
rect 42793 187584 42798 187640
rect 42854 187584 169708 187640
rect 42793 187582 169708 187584
rect 42793 187579 42859 187582
rect 169702 187580 169708 187582
rect 169772 187642 169778 187644
rect 170029 187642 170095 187645
rect 169772 187640 170095 187642
rect 169772 187584 170034 187640
rect 170090 187584 170095 187640
rect 169772 187582 170095 187584
rect 169772 187580 169778 187582
rect 170029 187579 170095 187582
rect 147070 187444 147076 187508
rect 147140 187506 147146 187508
rect 200113 187506 200179 187509
rect 147140 187504 200179 187506
rect 147140 187448 200118 187504
rect 200174 187448 200179 187504
rect 147140 187446 200179 187448
rect 147140 187444 147146 187446
rect 200113 187443 200179 187446
rect 214557 187506 214623 187509
rect 566641 187506 566707 187509
rect 214557 187504 566707 187506
rect 214557 187448 214562 187504
rect 214618 187448 566646 187504
rect 566702 187448 566707 187504
rect 214557 187446 566707 187448
rect 214557 187443 214623 187446
rect 566641 187443 566707 187446
rect 122966 187308 122972 187372
rect 123036 187370 123042 187372
rect 151169 187370 151235 187373
rect 123036 187368 151235 187370
rect 123036 187312 151174 187368
rect 151230 187312 151235 187368
rect 123036 187310 151235 187312
rect 123036 187308 123042 187310
rect 151169 187307 151235 187310
rect 174670 187308 174676 187372
rect 174740 187370 174746 187372
rect 207606 187370 207612 187372
rect 174740 187310 207612 187370
rect 174740 187308 174746 187310
rect 207606 187308 207612 187310
rect 207676 187370 207682 187372
rect 566457 187370 566523 187373
rect 207676 187368 566523 187370
rect 207676 187312 566462 187368
rect 566518 187312 566523 187368
rect 207676 187310 566523 187312
rect 207676 187308 207682 187310
rect 566457 187307 566523 187310
rect 113950 187172 113956 187236
rect 114020 187234 114026 187236
rect 147213 187234 147279 187237
rect 114020 187232 147279 187234
rect 114020 187176 147218 187232
rect 147274 187176 147279 187232
rect 114020 187174 147279 187176
rect 114020 187172 114026 187174
rect 147213 187171 147279 187174
rect 174854 187172 174860 187236
rect 174924 187234 174930 187236
rect 207473 187234 207539 187237
rect 572161 187234 572227 187237
rect 174924 187232 572227 187234
rect 174924 187176 207478 187232
rect 207534 187176 572166 187232
rect 572222 187176 572227 187232
rect 174924 187174 572227 187176
rect 174924 187172 174930 187174
rect 207473 187171 207539 187174
rect 572161 187171 572227 187174
rect 108430 187036 108436 187100
rect 108500 187098 108506 187100
rect 142981 187098 143047 187101
rect 108500 187096 143047 187098
rect 108500 187040 142986 187096
rect 143042 187040 143047 187096
rect 108500 187038 143047 187040
rect 108500 187036 108506 187038
rect 142981 187035 143047 187038
rect 168230 187036 168236 187100
rect 168300 187098 168306 187100
rect 201493 187098 201559 187101
rect 575013 187098 575079 187101
rect 168300 187096 575079 187098
rect 168300 187040 201498 187096
rect 201554 187040 575018 187096
rect 575074 187040 575079 187096
rect 168300 187038 575079 187040
rect 168300 187036 168306 187038
rect 201493 187035 201559 187038
rect 575013 187035 575079 187038
rect 112478 186900 112484 186964
rect 112548 186962 112554 186964
rect 147070 186962 147076 186964
rect 112548 186902 147076 186962
rect 112548 186900 112554 186902
rect 147070 186900 147076 186902
rect 147140 186900 147146 186964
rect 153469 186962 153535 186965
rect 187918 186962 187924 186964
rect 153469 186960 187924 186962
rect 153469 186904 153474 186960
rect 153530 186904 187924 186960
rect 153469 186902 187924 186904
rect 153469 186899 153535 186902
rect 187918 186900 187924 186902
rect 187988 186962 187994 186964
rect 569309 186962 569375 186965
rect 187988 186960 569375 186962
rect 187988 186904 569314 186960
rect 569370 186904 569375 186960
rect 187988 186902 569375 186904
rect 187988 186900 187994 186902
rect 569309 186899 569375 186902
rect 169334 186764 169340 186828
rect 169404 186826 169410 186828
rect 214557 186826 214623 186829
rect 169404 186824 214623 186826
rect 169404 186768 214562 186824
rect 214618 186768 214623 186824
rect 169404 186766 214623 186768
rect 169404 186764 169410 186766
rect 214557 186763 214623 186766
rect 144126 186220 144132 186284
rect 144196 186282 144202 186284
rect 144729 186282 144795 186285
rect 144196 186280 144795 186282
rect 144196 186224 144734 186280
rect 144790 186224 144795 186280
rect 144196 186222 144795 186224
rect 144196 186220 144202 186222
rect 144729 186219 144795 186222
rect 146886 186220 146892 186284
rect 146956 186282 146962 186284
rect 282913 186282 282979 186285
rect 146956 186280 282979 186282
rect 146956 186224 282918 186280
rect 282974 186224 282979 186280
rect 146956 186222 282979 186224
rect 146956 186220 146962 186222
rect 282913 186219 282979 186222
rect 49693 186146 49759 186149
rect 175222 186146 175228 186148
rect 49693 186144 175228 186146
rect 49693 186088 49698 186144
rect 49754 186088 175228 186144
rect 49693 186086 175228 186088
rect 49693 186083 49759 186086
rect 175222 186084 175228 186086
rect 175292 186146 175298 186148
rect 175641 186146 175707 186149
rect 175292 186144 175707 186146
rect 175292 186088 175646 186144
rect 175702 186088 175707 186144
rect 175292 186086 175707 186088
rect 175292 186084 175298 186086
rect 175641 186083 175707 186086
rect 168741 186010 168807 186013
rect 169150 186010 169156 186012
rect 168741 186008 169156 186010
rect 168741 185952 168746 186008
rect 168802 185952 169156 186008
rect 168741 185950 169156 185952
rect 168741 185947 168807 185950
rect 169150 185948 169156 185950
rect 169220 185948 169226 186012
rect 173750 185812 173756 185876
rect 173820 185874 173826 185876
rect 217041 185874 217107 185877
rect 567929 185874 567995 185877
rect 173820 185872 567995 185874
rect 173820 185816 217046 185872
rect 217102 185816 567934 185872
rect 567990 185816 567995 185872
rect 173820 185814 567995 185816
rect 173820 185812 173826 185814
rect 217041 185811 217107 185814
rect 567929 185811 567995 185814
rect 174486 185676 174492 185740
rect 174556 185738 174562 185740
rect 208669 185738 208735 185741
rect 570781 185738 570847 185741
rect 174556 185736 570847 185738
rect 174556 185680 208674 185736
rect 208730 185680 570786 185736
rect 570842 185680 570847 185736
rect 174556 185678 570847 185680
rect 174556 185676 174562 185678
rect 208669 185675 208735 185678
rect 570781 185675 570847 185678
rect 580257 185738 580323 185741
rect 583520 185738 584960 185828
rect 580257 185736 584960 185738
rect 580257 185680 580262 185736
rect 580318 185680 584960 185736
rect 580257 185678 584960 185680
rect 580257 185675 580323 185678
rect 112662 185540 112668 185604
rect 112732 185602 112738 185604
rect 146886 185602 146892 185604
rect 112732 185542 146892 185602
rect 112732 185540 112738 185542
rect 146886 185540 146892 185542
rect 146956 185540 146962 185604
rect 148910 185540 148916 185604
rect 148980 185602 148986 185604
rect 189206 185602 189212 185604
rect 148980 185542 189212 185602
rect 148980 185540 148986 185542
rect 189206 185540 189212 185542
rect 189276 185602 189282 185604
rect 580993 185602 581059 185605
rect 189276 185600 581059 185602
rect 189276 185544 580998 185600
rect 581054 185544 581059 185600
rect 583520 185588 584960 185678
rect 189276 185542 581059 185544
rect 189276 185540 189282 185542
rect 580993 185539 581059 185542
rect -960 185058 480 185148
rect 3417 185058 3483 185061
rect -960 185056 3483 185058
rect -960 185000 3422 185056
rect 3478 185000 3483 185056
rect -960 184998 3483 185000
rect -960 184908 480 184998
rect 3417 184995 3483 184998
rect 162710 184452 162716 184516
rect 162780 184514 162786 184516
rect 183369 184514 183435 184517
rect 444373 184514 444439 184517
rect 162780 184512 444439 184514
rect 162780 184456 183374 184512
rect 183430 184456 444378 184512
rect 444434 184456 444439 184512
rect 162780 184454 444439 184456
rect 162780 184452 162786 184454
rect 183369 184451 183435 184454
rect 444373 184451 444439 184454
rect 163998 184316 164004 184380
rect 164068 184378 164074 184380
rect 217317 184378 217383 184381
rect 561029 184378 561095 184381
rect 164068 184376 561095 184378
rect 164068 184320 217322 184376
rect 217378 184320 561034 184376
rect 561090 184320 561095 184376
rect 164068 184318 561095 184320
rect 164068 184316 164074 184318
rect 217317 184315 217383 184318
rect 561029 184315 561095 184318
rect 168966 184180 168972 184244
rect 169036 184242 169042 184244
rect 203558 184242 203564 184244
rect 169036 184182 203564 184242
rect 169036 184180 169042 184182
rect 203558 184180 203564 184182
rect 203628 184242 203634 184244
rect 552657 184242 552723 184245
rect 203628 184240 552723 184242
rect 203628 184184 552662 184240
rect 552718 184184 552723 184240
rect 203628 184182 552723 184184
rect 203628 184180 203634 184182
rect 552657 184179 552723 184182
rect 139025 183564 139091 183565
rect 138974 183562 138980 183564
rect 138934 183502 138980 183562
rect 139044 183560 139091 183564
rect 409873 183562 409939 183565
rect 139086 183504 139091 183560
rect 138974 183500 138980 183502
rect 139044 183500 139091 183504
rect 139025 183499 139091 183500
rect 142110 183560 409939 183562
rect 142110 183504 409878 183560
rect 409934 183504 409939 183560
rect 142110 183502 409939 183504
rect 107142 182820 107148 182884
rect 107212 182882 107218 182884
rect 139894 182882 139900 182884
rect 107212 182822 139900 182882
rect 107212 182820 107218 182822
rect 139894 182820 139900 182822
rect 139964 182882 139970 182884
rect 142110 182882 142170 183502
rect 409873 183499 409939 183502
rect 144177 183426 144243 183429
rect 144678 183426 144684 183428
rect 144177 183424 144684 183426
rect 144177 183368 144182 183424
rect 144238 183368 144684 183424
rect 144177 183366 144684 183368
rect 144177 183363 144243 183366
rect 144678 183364 144684 183366
rect 144748 183364 144754 183428
rect 217225 183426 217291 183429
rect 463693 183426 463759 183429
rect 200070 183424 463759 183426
rect 200070 183368 217230 183424
rect 217286 183368 463698 183424
rect 463754 183368 463759 183424
rect 200070 183366 463759 183368
rect 159030 183228 159036 183292
rect 159100 183290 159106 183292
rect 200070 183290 200130 183366
rect 217225 183363 217291 183366
rect 463693 183363 463759 183366
rect 218145 183290 218211 183293
rect 489913 183290 489979 183293
rect 159100 183230 200130 183290
rect 215710 183288 489979 183290
rect 215710 183232 218150 183288
rect 218206 183232 489918 183288
rect 489974 183232 489979 183288
rect 215710 183230 489979 183232
rect 159100 183228 159106 183230
rect 154062 183092 154068 183156
rect 154132 183154 154138 183156
rect 215710 183154 215770 183230
rect 218145 183227 218211 183230
rect 489913 183227 489979 183230
rect 154132 183094 215770 183154
rect 218237 183154 218303 183157
rect 582557 183154 582623 183157
rect 218237 183152 582623 183154
rect 218237 183096 218242 183152
rect 218298 183096 582562 183152
rect 582618 183096 582623 183152
rect 218237 183094 582623 183096
rect 154132 183092 154138 183094
rect 218237 183091 218303 183094
rect 582557 183091 582623 183094
rect 158897 183018 158963 183021
rect 185710 183018 185716 183020
rect 158897 183016 185716 183018
rect 158897 182960 158902 183016
rect 158958 182960 185716 183016
rect 158897 182958 185716 182960
rect 158897 182955 158963 182958
rect 185710 182956 185716 182958
rect 185780 183018 185786 183020
rect 565077 183018 565143 183021
rect 185780 183016 565143 183018
rect 185780 182960 565082 183016
rect 565138 182960 565143 183016
rect 185780 182958 565143 182960
rect 185780 182956 185786 182958
rect 565077 182955 565143 182958
rect 139964 182822 142170 182882
rect 139964 182820 139970 182822
rect 154246 182820 154252 182884
rect 154316 182882 154322 182884
rect 186078 182882 186084 182884
rect 154316 182822 186084 182882
rect 154316 182820 154322 182822
rect 186078 182820 186084 182822
rect 186148 182882 186154 182884
rect 582465 182882 582531 182885
rect 186148 182880 582531 182882
rect 186148 182824 582470 182880
rect 582526 182824 582531 182880
rect 186148 182822 582531 182824
rect 186148 182820 186154 182822
rect 582465 182819 582531 182822
rect 144177 182746 144243 182749
rect 309133 182746 309199 182749
rect 144177 182744 309199 182746
rect 144177 182688 144182 182744
rect 144238 182688 309138 182744
rect 309194 182688 309199 182744
rect 144177 182686 309199 182688
rect 144177 182683 144243 182686
rect 309133 182683 309199 182686
rect 157190 182548 157196 182612
rect 157260 182610 157266 182612
rect 218237 182610 218303 182613
rect 157260 182608 218303 182610
rect 157260 182552 218242 182608
rect 218298 182552 218303 182608
rect 157260 182550 218303 182552
rect 157260 182548 157266 182550
rect 218237 182547 218303 182550
rect 108614 182140 108620 182204
rect 108684 182202 108690 182204
rect 143441 182202 143507 182205
rect 108684 182200 143507 182202
rect 108684 182144 143446 182200
rect 143502 182144 143507 182200
rect 108684 182142 143507 182144
rect 108684 182140 108690 182142
rect 143441 182139 143507 182142
rect 149697 182066 149763 182069
rect 150014 182066 150020 182068
rect 149697 182064 150020 182066
rect 149697 182008 149702 182064
rect 149758 182008 150020 182064
rect 149697 182006 150020 182008
rect 149697 182003 149763 182006
rect 150014 182004 150020 182006
rect 150084 182066 150090 182068
rect 459553 182066 459619 182069
rect 150084 182064 459619 182066
rect 150084 182008 459558 182064
rect 459614 182008 459619 182064
rect 150084 182006 459619 182008
rect 150084 182004 150090 182006
rect 459553 182003 459619 182006
rect 580165 181658 580231 181661
rect 583520 181658 584960 181748
rect 580165 181656 584960 181658
rect 580165 181600 580170 181656
rect 580226 181600 584960 181656
rect 580165 181598 584960 181600
rect 580165 181595 580231 181598
rect 583520 181508 584960 181598
rect 151670 181324 151676 181388
rect 151740 181386 151746 181388
rect 216857 181386 216923 181389
rect 539593 181386 539659 181389
rect 151740 181384 539659 181386
rect 151740 181328 216862 181384
rect 216918 181328 539598 181384
rect 539654 181328 539659 181384
rect 151740 181326 539659 181328
rect 151740 181324 151746 181326
rect 216857 181323 216923 181326
rect 539593 181323 539659 181326
rect -960 180978 480 181068
rect 3417 180978 3483 180981
rect -960 180976 3483 180978
rect -960 180920 3422 180976
rect 3478 180920 3483 180976
rect -960 180918 3483 180920
rect -960 180828 480 180918
rect 3417 180915 3483 180918
rect 100518 180916 100524 180980
rect 100588 180978 100594 180980
rect 120717 180978 120783 180981
rect 100588 180976 120783 180978
rect 100588 180920 120722 180976
rect 120778 180920 120783 180976
rect 100588 180918 120783 180920
rect 100588 180916 100594 180918
rect 120717 180915 120783 180918
rect 104566 180780 104572 180844
rect 104636 180842 104642 180844
rect 138790 180842 138796 180844
rect 104636 180782 138796 180842
rect 104636 180780 104642 180782
rect 138790 180780 138796 180782
rect 138860 180780 138866 180844
rect 137870 180644 137876 180708
rect 137940 180706 137946 180708
rect 582925 180706 582991 180709
rect 137940 180704 582991 180706
rect 137940 180648 582930 180704
rect 582986 180648 582991 180704
rect 137940 180646 582991 180648
rect 137940 180644 137946 180646
rect 582925 180643 582991 180646
rect 142521 180570 142587 180573
rect 565169 180570 565235 180573
rect 142521 180568 565235 180570
rect 142521 180512 142526 180568
rect 142582 180512 565174 180568
rect 565230 180512 565235 180568
rect 142521 180510 565235 180512
rect 142521 180507 142587 180510
rect 565169 180507 565235 180510
rect 138790 180372 138796 180436
rect 138860 180434 138866 180436
rect 494697 180434 494763 180437
rect 138860 180432 494763 180434
rect 138860 180376 494702 180432
rect 494758 180376 494763 180432
rect 138860 180374 494763 180376
rect 138860 180372 138866 180374
rect 494697 180371 494763 180374
rect 481633 180298 481699 180301
rect 142110 180296 481699 180298
rect 142110 180240 481638 180296
rect 481694 180240 481699 180296
rect 142110 180238 481699 180240
rect 104750 180100 104756 180164
rect 104820 180162 104826 180164
rect 138606 180162 138612 180164
rect 104820 180102 138612 180162
rect 104820 180100 104826 180102
rect 138606 180100 138612 180102
rect 138676 180162 138682 180164
rect 142110 180162 142170 180238
rect 481633 180235 481699 180238
rect 138676 180102 142170 180162
rect 138676 180100 138682 180102
rect 107326 179964 107332 180028
rect 107396 180026 107402 180028
rect 142521 180026 142587 180029
rect 107396 180024 142587 180026
rect 107396 179968 142526 180024
rect 142582 179968 142587 180024
rect 107396 179966 142587 179968
rect 107396 179964 107402 179966
rect 142521 179963 142587 179966
rect 106038 179692 106044 179756
rect 106108 179754 106114 179756
rect 127709 179754 127775 179757
rect 106108 179752 127775 179754
rect 106108 179696 127714 179752
rect 127770 179696 127775 179752
rect 106108 179694 127775 179696
rect 106108 179692 106114 179694
rect 127709 179691 127775 179694
rect 103278 179556 103284 179620
rect 103348 179618 103354 179620
rect 124765 179618 124831 179621
rect 103348 179616 124831 179618
rect 103348 179560 124770 179616
rect 124826 179560 124831 179616
rect 103348 179558 124831 179560
rect 103348 179556 103354 179558
rect 124765 179555 124831 179558
rect 99046 179420 99052 179484
rect 99116 179482 99122 179484
rect 123477 179482 123543 179485
rect 124029 179482 124095 179485
rect 99116 179480 124095 179482
rect 99116 179424 123482 179480
rect 123538 179424 124034 179480
rect 124090 179424 124095 179480
rect 99116 179422 124095 179424
rect 99116 179420 99122 179422
rect 123477 179419 123543 179422
rect 124029 179419 124095 179422
rect 136214 179420 136220 179484
rect 136284 179482 136290 179484
rect 136541 179482 136607 179485
rect 136284 179480 136607 179482
rect 136284 179424 136546 179480
rect 136602 179424 136607 179480
rect 136284 179422 136607 179424
rect 136284 179420 136290 179422
rect 136541 179419 136607 179422
rect 137277 179482 137343 179485
rect 137870 179482 137876 179484
rect 137277 179480 137876 179482
rect 137277 179424 137282 179480
rect 137338 179424 137876 179480
rect 137277 179422 137876 179424
rect 137277 179419 137343 179422
rect 137870 179420 137876 179422
rect 137940 179420 137946 179484
rect 166206 178876 166212 178940
rect 166276 178938 166282 178940
rect 214189 178938 214255 178941
rect 570689 178938 570755 178941
rect 166276 178936 570755 178938
rect 166276 178880 214194 178936
rect 214250 178880 570694 178936
rect 570750 178880 570755 178936
rect 166276 178878 570755 178880
rect 166276 178876 166282 178878
rect 214189 178875 214255 178878
rect 570689 178875 570755 178878
rect 171726 178740 171732 178804
rect 171796 178802 171802 178804
rect 203006 178802 203012 178804
rect 171796 178742 203012 178802
rect 171796 178740 171802 178742
rect 203006 178740 203012 178742
rect 203076 178802 203082 178804
rect 573357 178802 573423 178805
rect 203076 178800 573423 178802
rect 203076 178744 573362 178800
rect 573418 178744 573423 178800
rect 203076 178742 573423 178744
rect 203076 178740 203082 178742
rect 573357 178739 573423 178742
rect 165102 178604 165108 178668
rect 165172 178666 165178 178668
rect 176561 178666 176627 178669
rect 556889 178666 556955 178669
rect 165172 178664 556955 178666
rect 165172 178608 176566 178664
rect 176622 178608 556894 178664
rect 556950 178608 556955 178664
rect 165172 178606 556955 178608
rect 165172 178604 165178 178606
rect 176561 178603 176627 178606
rect 556889 178603 556955 178606
rect 140998 177924 141004 177988
rect 141068 177986 141074 177988
rect 141417 177986 141483 177989
rect 544469 177986 544535 177989
rect 141068 177984 544535 177986
rect 141068 177928 141422 177984
rect 141478 177928 544474 177984
rect 544530 177928 544535 177984
rect 141068 177926 544535 177928
rect 141068 177924 141074 177926
rect 141417 177923 141483 177926
rect 544469 177923 544535 177926
rect 136030 177788 136036 177852
rect 136100 177850 136106 177852
rect 136449 177850 136515 177853
rect 136100 177848 136515 177850
rect 136100 177792 136454 177848
rect 136510 177792 136515 177848
rect 136100 177790 136515 177792
rect 136100 177788 136106 177790
rect 136449 177787 136515 177790
rect -960 177578 480 177668
rect 3325 177578 3391 177581
rect -960 177576 3391 177578
rect -960 177520 3330 177576
rect 3386 177520 3391 177576
rect -960 177518 3391 177520
rect -960 177428 480 177518
rect 3325 177515 3391 177518
rect 580165 177578 580231 177581
rect 583520 177578 584960 177668
rect 580165 177576 584960 177578
rect 580165 177520 580170 177576
rect 580226 177520 584960 177576
rect 580165 177518 584960 177520
rect 580165 177515 580231 177518
rect 583520 177428 584960 177518
rect 122230 176564 122236 176628
rect 122300 176626 122306 176628
rect 548517 176626 548583 176629
rect 122300 176624 548583 176626
rect 122300 176568 548522 176624
rect 548578 176568 548583 176624
rect 122300 176566 548583 176568
rect 122300 176564 122306 176566
rect 548517 176563 548583 176566
rect 121126 176428 121132 176492
rect 121196 176490 121202 176492
rect 140957 176490 141023 176493
rect 558269 176490 558335 176493
rect 121196 176488 558335 176490
rect 121196 176432 140962 176488
rect 141018 176432 558274 176488
rect 558330 176432 558335 176488
rect 121196 176430 558335 176432
rect 121196 176428 121202 176430
rect 140957 176427 141023 176430
rect 558269 176427 558335 176430
rect 102910 176292 102916 176356
rect 102980 176354 102986 176356
rect 137134 176354 137140 176356
rect 102980 176294 137140 176354
rect 102980 176292 102986 176294
rect 137134 176292 137140 176294
rect 137204 176354 137210 176356
rect 544377 176354 544443 176357
rect 137204 176352 544443 176354
rect 137204 176296 544382 176352
rect 544438 176296 544443 176352
rect 137204 176294 544443 176296
rect 137204 176292 137210 176294
rect 544377 176291 544443 176294
rect 103094 176156 103100 176220
rect 103164 176218 103170 176220
rect 136817 176218 136883 176221
rect 382273 176218 382339 176221
rect 103164 176216 382339 176218
rect 103164 176160 136822 176216
rect 136878 176160 382278 176216
rect 382334 176160 382339 176216
rect 103164 176158 382339 176160
rect 103164 176156 103170 176158
rect 136817 176155 136883 176158
rect 382273 176155 382339 176158
rect 124806 176020 124812 176084
rect 124876 176082 124882 176084
rect 140865 176082 140931 176085
rect 367093 176082 367159 176085
rect 124876 176080 367159 176082
rect 124876 176024 140870 176080
rect 140926 176024 367098 176080
rect 367154 176024 367159 176080
rect 124876 176022 367159 176024
rect 124876 176020 124882 176022
rect 140865 176019 140931 176022
rect 367093 176019 367159 176022
rect 121310 175884 121316 175948
rect 121380 175946 121386 175948
rect 135846 175946 135852 175948
rect 121380 175886 135852 175946
rect 121380 175884 121386 175886
rect 135846 175884 135852 175886
rect 135916 175946 135922 175948
rect 351913 175946 351979 175949
rect 135916 175944 351979 175946
rect 135916 175888 351918 175944
rect 351974 175888 351979 175944
rect 135916 175886 351979 175888
rect 135916 175884 135922 175886
rect 351913 175883 351979 175886
rect -960 173498 480 173588
rect 3417 173498 3483 173501
rect -960 173496 3483 173498
rect -960 173440 3422 173496
rect 3478 173440 3483 173496
rect -960 173438 3483 173440
rect -960 173348 480 173438
rect 3417 173435 3483 173438
rect 580165 173498 580231 173501
rect 583520 173498 584960 173588
rect 580165 173496 584960 173498
rect 580165 173440 580170 173496
rect 580226 173440 584960 173496
rect 580165 173438 584960 173440
rect 580165 173435 580231 173438
rect 583520 173348 584960 173438
rect -960 169418 480 169508
rect 3141 169418 3207 169421
rect -960 169416 3207 169418
rect -960 169360 3146 169416
rect 3202 169360 3207 169416
rect -960 169358 3207 169360
rect -960 169268 480 169358
rect 3141 169355 3207 169358
rect 580257 169418 580323 169421
rect 583520 169418 584960 169508
rect 580257 169416 584960 169418
rect 580257 169360 580262 169416
rect 580318 169360 584960 169416
rect 580257 169358 584960 169360
rect 580257 169355 580323 169358
rect 583520 169268 584960 169358
rect -960 165338 480 165428
rect 2773 165338 2839 165341
rect -960 165336 2839 165338
rect -960 165280 2778 165336
rect 2834 165280 2839 165336
rect -960 165278 2839 165280
rect -960 165188 480 165278
rect 2773 165275 2839 165278
rect 580165 165338 580231 165341
rect 583520 165338 584960 165428
rect 580165 165336 584960 165338
rect 580165 165280 580170 165336
rect 580226 165280 584960 165336
rect 580165 165278 584960 165280
rect 580165 165275 580231 165278
rect 583520 165188 584960 165278
rect 580165 161938 580231 161941
rect 583520 161938 584960 162028
rect 580165 161936 584960 161938
rect 580165 161880 580170 161936
rect 580226 161880 584960 161936
rect 580165 161878 584960 161880
rect 580165 161875 580231 161878
rect 583520 161788 584960 161878
rect -960 161258 480 161348
rect 3509 161258 3575 161261
rect -960 161256 3575 161258
rect -960 161200 3514 161256
rect 3570 161200 3575 161256
rect -960 161198 3575 161200
rect -960 161108 480 161198
rect 3509 161195 3575 161198
rect 583520 157708 584960 157948
rect -960 157178 480 157268
rect 3509 157178 3575 157181
rect -960 157176 3575 157178
rect -960 157120 3514 157176
rect 3570 157120 3575 157176
rect -960 157118 3575 157120
rect -960 157028 480 157118
rect 3509 157115 3575 157118
rect 579613 153778 579679 153781
rect 583520 153778 584960 153868
rect 579613 153776 584960 153778
rect 579613 153720 579618 153776
rect 579674 153720 584960 153776
rect 579613 153718 584960 153720
rect 579613 153715 579679 153718
rect 583520 153628 584960 153718
rect -960 153098 480 153188
rect 3509 153098 3575 153101
rect -960 153096 3575 153098
rect -960 153040 3514 153096
rect 3570 153040 3575 153096
rect -960 153038 3575 153040
rect -960 152948 480 153038
rect 3509 153035 3575 153038
rect 580165 149698 580231 149701
rect 583520 149698 584960 149788
rect 580165 149696 584960 149698
rect 580165 149640 580170 149696
rect 580226 149640 584960 149696
rect 580165 149638 584960 149640
rect 580165 149635 580231 149638
rect 583520 149548 584960 149638
rect -960 149018 480 149108
rect 3417 149018 3483 149021
rect -960 149016 3483 149018
rect -960 148960 3422 149016
rect 3478 148960 3483 149016
rect -960 148958 3483 148960
rect -960 148868 480 148958
rect 3417 148955 3483 148958
rect 100334 148548 100340 148612
rect 100404 148610 100410 148612
rect 126973 148610 127039 148613
rect 100404 148608 127039 148610
rect 100404 148552 126978 148608
rect 127034 148552 127039 148608
rect 100404 148550 127039 148552
rect 100404 148548 100410 148550
rect 126973 148547 127039 148550
rect 111006 148412 111012 148476
rect 111076 148474 111082 148476
rect 142797 148474 142863 148477
rect 111076 148472 142863 148474
rect 111076 148416 142802 148472
rect 142858 148416 142863 148472
rect 111076 148414 142863 148416
rect 111076 148412 111082 148414
rect 142797 148411 142863 148414
rect 168465 148474 168531 148477
rect 203517 148474 203583 148477
rect 168465 148472 203583 148474
rect 168465 148416 168470 148472
rect 168526 148416 203522 148472
rect 203578 148416 203583 148472
rect 168465 148414 203583 148416
rect 168465 148411 168531 148414
rect 203517 148411 203583 148414
rect 106958 148276 106964 148340
rect 107028 148338 107034 148340
rect 148133 148338 148199 148341
rect 107028 148336 148199 148338
rect 107028 148280 148138 148336
rect 148194 148280 148199 148336
rect 107028 148278 148199 148280
rect 107028 148276 107034 148278
rect 148133 148275 148199 148278
rect 152549 148338 152615 148341
rect 216121 148338 216187 148341
rect 152549 148336 216187 148338
rect 152549 148280 152554 148336
rect 152610 148280 216126 148336
rect 216182 148280 216187 148336
rect 152549 148278 216187 148280
rect 152549 148275 152615 148278
rect 216121 148275 216187 148278
rect 146293 147794 146359 147797
rect 580533 147794 580599 147797
rect 146293 147792 580599 147794
rect 146293 147736 146298 147792
rect 146354 147736 580538 147792
rect 580594 147736 580599 147792
rect 146293 147734 580599 147736
rect 146293 147731 146359 147734
rect 580533 147731 580599 147734
rect 176561 146978 176627 146981
rect 198958 146978 198964 146980
rect 176561 146976 198964 146978
rect 176561 146920 176566 146976
rect 176622 146920 198964 146976
rect 176561 146918 198964 146920
rect 176561 146915 176627 146918
rect 198958 146916 198964 146918
rect 199028 146916 199034 146980
rect 111558 145964 111564 146028
rect 111628 146026 111634 146028
rect 130101 146026 130167 146029
rect 111628 146024 130167 146026
rect 111628 145968 130106 146024
rect 130162 145968 130167 146024
rect 111628 145966 130167 145968
rect 111628 145964 111634 145966
rect 130101 145963 130167 145966
rect 182265 146026 182331 146029
rect 197486 146026 197492 146028
rect 182265 146024 197492 146026
rect 182265 145968 182270 146024
rect 182326 145968 197492 146024
rect 182265 145966 197492 145968
rect 182265 145963 182331 145966
rect 197486 145964 197492 145966
rect 197556 145964 197562 146028
rect 111374 145828 111380 145892
rect 111444 145890 111450 145892
rect 132585 145890 132651 145893
rect 111444 145888 132651 145890
rect 111444 145832 132590 145888
rect 132646 145832 132651 145888
rect 111444 145830 132651 145832
rect 111444 145828 111450 145830
rect 132585 145827 132651 145830
rect 171501 145890 171567 145893
rect 195329 145890 195395 145893
rect 171501 145888 195395 145890
rect 171501 145832 171506 145888
rect 171562 145832 195334 145888
rect 195390 145832 195395 145888
rect 171501 145830 195395 145832
rect 171501 145827 171567 145830
rect 195329 145827 195395 145830
rect 112846 145692 112852 145756
rect 112916 145754 112922 145756
rect 136725 145754 136791 145757
rect 112916 145752 136791 145754
rect 112916 145696 136730 145752
rect 136786 145696 136791 145752
rect 112916 145694 136791 145696
rect 112916 145692 112922 145694
rect 136725 145691 136791 145694
rect 169017 145754 169083 145757
rect 196198 145754 196204 145756
rect 169017 145752 196204 145754
rect 169017 145696 169022 145752
rect 169078 145696 196204 145752
rect 169017 145694 196204 145696
rect 169017 145691 169083 145694
rect 196198 145692 196204 145694
rect 196268 145692 196274 145756
rect 116577 145618 116643 145621
rect 150065 145618 150131 145621
rect 116577 145616 150131 145618
rect 116577 145560 116582 145616
rect 116638 145560 150070 145616
rect 150126 145560 150131 145616
rect 116577 145558 150131 145560
rect 116577 145555 116643 145558
rect 150065 145555 150131 145558
rect 164417 145618 164483 145621
rect 196985 145618 197051 145621
rect 164417 145616 197051 145618
rect 164417 145560 164422 145616
rect 164478 145560 196990 145616
rect 197046 145560 197051 145616
rect 164417 145558 197051 145560
rect 164417 145555 164483 145558
rect 196985 145555 197051 145558
rect 580165 145618 580231 145621
rect 583520 145618 584960 145708
rect 580165 145616 584960 145618
rect 580165 145560 580170 145616
rect 580226 145560 584960 145616
rect 580165 145558 584960 145560
rect 580165 145555 580231 145558
rect 583520 145468 584960 145558
rect -960 144938 480 145028
rect 3417 144938 3483 144941
rect -960 144936 3483 144938
rect -960 144880 3422 144936
rect 3478 144880 3483 144936
rect -960 144878 3483 144880
rect -960 144788 480 144878
rect 3417 144875 3483 144878
rect 111558 144332 111564 144396
rect 111628 144394 111634 144396
rect 144177 144394 144243 144397
rect 111628 144392 144243 144394
rect 111628 144336 144182 144392
rect 144238 144336 144243 144392
rect 111628 144334 144243 144336
rect 111628 144332 111634 144334
rect 144177 144331 144243 144334
rect 184749 144394 184815 144397
rect 196566 144394 196572 144396
rect 184749 144392 196572 144394
rect 184749 144336 184754 144392
rect 184810 144336 196572 144392
rect 184749 144334 196572 144336
rect 184749 144331 184815 144334
rect 196566 144332 196572 144334
rect 196636 144332 196642 144396
rect 116526 144196 116532 144260
rect 116596 144258 116602 144260
rect 149697 144258 149763 144261
rect 116596 144256 149763 144258
rect 116596 144200 149702 144256
rect 149758 144200 149763 144256
rect 116596 144198 149763 144200
rect 116596 144196 116602 144198
rect 149697 144195 149763 144198
rect 161974 144196 161980 144260
rect 162044 144258 162050 144260
rect 187509 144258 187575 144261
rect 162044 144256 187575 144258
rect 162044 144200 187514 144256
rect 187570 144200 187575 144256
rect 162044 144198 187575 144200
rect 162044 144196 162050 144198
rect 187509 144195 187575 144198
rect 113766 144060 113772 144124
rect 113836 144122 113842 144124
rect 149513 144122 149579 144125
rect 113836 144120 149579 144122
rect 113836 144064 149518 144120
rect 149574 144064 149579 144120
rect 113836 144062 149579 144064
rect 113836 144060 113842 144062
rect 149513 144059 149579 144062
rect 157977 144122 158043 144125
rect 192150 144122 192156 144124
rect 157977 144120 192156 144122
rect 157977 144064 157982 144120
rect 158038 144064 192156 144120
rect 157977 144062 192156 144064
rect 157977 144059 158043 144062
rect 192150 144060 192156 144062
rect 192220 144060 192226 144124
rect 169753 143578 169819 143581
rect 192385 143578 192451 143581
rect 192845 143578 192911 143581
rect 169753 143576 192911 143578
rect 169753 143520 169758 143576
rect 169814 143520 192390 143576
rect 192446 143520 192850 143576
rect 192906 143520 192911 143576
rect 169753 143518 192911 143520
rect 169753 143515 169819 143518
rect 192385 143515 192451 143518
rect 192845 143515 192911 143518
rect 178585 143442 178651 143445
rect 186773 143442 186839 143445
rect 178585 143440 186839 143442
rect 178585 143384 178590 143440
rect 178646 143384 186778 143440
rect 186834 143384 186839 143440
rect 178585 143382 186839 143384
rect 178585 143379 178651 143382
rect 186773 143379 186839 143382
rect 186957 143442 187023 143445
rect 187182 143442 187188 143444
rect 186957 143440 187188 143442
rect 186957 143384 186962 143440
rect 187018 143384 187188 143440
rect 186957 143382 187188 143384
rect 186957 143379 187023 143382
rect 187182 143380 187188 143382
rect 187252 143380 187258 143444
rect 196014 143306 196020 143308
rect 186270 143246 196020 143306
rect 186270 143173 186330 143246
rect 196014 143244 196020 143246
rect 196084 143244 196090 143308
rect 114001 143170 114067 143173
rect 124397 143170 124463 143173
rect 114001 143168 124463 143170
rect 114001 143112 114006 143168
rect 114062 143112 124402 143168
rect 124458 143112 124463 143168
rect 114001 143110 124463 143112
rect 114001 143107 114067 143110
rect 124397 143107 124463 143110
rect 186221 143168 186330 143173
rect 186221 143112 186226 143168
rect 186282 143112 186330 143168
rect 186221 143110 186330 143112
rect 186221 143107 186287 143110
rect 186998 143108 187004 143172
rect 187068 143170 187074 143172
rect 187601 143170 187667 143173
rect 187068 143168 187667 143170
rect 187068 143112 187606 143168
rect 187662 143112 187667 143168
rect 187068 143110 187667 143112
rect 187068 143108 187074 143110
rect 187601 143107 187667 143110
rect 116894 142972 116900 143036
rect 116964 143034 116970 143036
rect 135989 143034 136055 143037
rect 116964 143032 136055 143034
rect 116964 142976 135994 143032
rect 136050 142976 136055 143032
rect 116964 142974 136055 142976
rect 116964 142972 116970 142974
rect 135989 142971 136055 142974
rect 179413 143034 179479 143037
rect 186589 143034 186655 143037
rect 179413 143032 186655 143034
rect 179413 142976 179418 143032
rect 179474 142976 186594 143032
rect 186650 142976 186655 143032
rect 179413 142974 186655 142976
rect 179413 142971 179479 142974
rect 186589 142971 186655 142974
rect 186773 143034 186839 143037
rect 192109 143034 192175 143037
rect 186773 143032 192175 143034
rect 186773 142976 186778 143032
rect 186834 142976 192114 143032
rect 192170 142976 192175 143032
rect 186773 142974 192175 142976
rect 186773 142971 186839 142974
rect 192109 142971 192175 142974
rect 118550 142836 118556 142900
rect 118620 142898 118626 142900
rect 148409 142898 148475 142901
rect 118620 142896 148475 142898
rect 118620 142840 148414 142896
rect 148470 142840 148475 142896
rect 118620 142838 148475 142840
rect 118620 142836 118626 142838
rect 148409 142835 148475 142838
rect 178861 142898 178927 142901
rect 193254 142898 193260 142900
rect 178861 142896 193260 142898
rect 178861 142840 178866 142896
rect 178922 142840 193260 142896
rect 178861 142838 193260 142840
rect 178861 142835 178927 142838
rect 193254 142836 193260 142838
rect 193324 142836 193330 142900
rect 115381 142762 115447 142765
rect 146753 142762 146819 142765
rect 115381 142760 146819 142762
rect 115381 142704 115386 142760
rect 115442 142704 146758 142760
rect 146814 142704 146819 142760
rect 115381 142702 146819 142704
rect 115381 142699 115447 142702
rect 146753 142699 146819 142702
rect 183461 142762 183527 142765
rect 191782 142762 191788 142764
rect 183461 142760 191788 142762
rect 183461 142704 183466 142760
rect 183522 142704 191788 142760
rect 183461 142702 191788 142704
rect 183461 142699 183527 142702
rect 191782 142700 191788 142702
rect 191852 142762 191858 142764
rect 579613 142762 579679 142765
rect 191852 142760 579679 142762
rect 191852 142704 579618 142760
rect 579674 142704 579679 142760
rect 191852 142702 579679 142704
rect 191852 142700 191858 142702
rect 579613 142699 579679 142702
rect 184657 142626 184723 142629
rect 195421 142626 195487 142629
rect 184657 142624 195487 142626
rect 184657 142568 184662 142624
rect 184718 142568 195426 142624
rect 195482 142568 195487 142624
rect 184657 142566 195487 142568
rect 184657 142563 184723 142566
rect 195421 142563 195487 142566
rect 186589 142490 186655 142493
rect 193581 142490 193647 142493
rect 186589 142488 193647 142490
rect 186589 142432 186594 142488
rect 186650 142432 193586 142488
rect 193642 142432 193647 142488
rect 186589 142430 193647 142432
rect 186589 142427 186655 142430
rect 193581 142427 193647 142430
rect 157241 142354 157307 142357
rect 190453 142354 190519 142357
rect 157241 142352 190519 142354
rect 157241 142296 157246 142352
rect 157302 142296 190458 142352
rect 190514 142296 190519 142352
rect 157241 142294 190519 142296
rect 157241 142291 157307 142294
rect 190453 142291 190519 142294
rect 112846 141884 112852 141948
rect 112916 141946 112922 141948
rect 130837 141946 130903 141949
rect 112916 141944 130903 141946
rect 112916 141888 130842 141944
rect 130898 141888 130903 141944
rect 112916 141886 130903 141888
rect 112916 141884 112922 141886
rect 130837 141883 130903 141886
rect 181989 141946 182055 141949
rect 192661 141946 192727 141949
rect 181989 141944 192727 141946
rect 181989 141888 181994 141944
rect 182050 141888 192666 141944
rect 192722 141888 192727 141944
rect 181989 141886 192727 141888
rect 181989 141883 182055 141886
rect 192661 141883 192727 141886
rect 97073 141810 97139 141813
rect 134517 141810 134583 141813
rect 97073 141808 134583 141810
rect 97073 141752 97078 141808
rect 97134 141752 134522 141808
rect 134578 141752 134583 141808
rect 97073 141750 134583 141752
rect 97073 141747 97139 141750
rect 134517 141747 134583 141750
rect 165613 141810 165679 141813
rect 207749 141810 207815 141813
rect 165613 141808 207815 141810
rect 165613 141752 165618 141808
rect 165674 141752 207754 141808
rect 207810 141752 207815 141808
rect 165613 141750 207815 141752
rect 165613 141747 165679 141750
rect 207749 141747 207815 141750
rect 118550 141612 118556 141676
rect 118620 141674 118626 141676
rect 178033 141674 178099 141677
rect 118620 141672 178099 141674
rect 118620 141616 178038 141672
rect 178094 141616 178099 141672
rect 118620 141614 178099 141616
rect 118620 141612 118626 141614
rect 178033 141611 178099 141614
rect 181897 141674 181963 141677
rect 193438 141674 193444 141676
rect 181897 141672 193444 141674
rect 181897 141616 181902 141672
rect 181958 141616 193444 141672
rect 181897 141614 193444 141616
rect 181897 141611 181963 141614
rect 193438 141612 193444 141614
rect 193508 141612 193514 141676
rect 118182 141476 118188 141540
rect 118252 141538 118258 141540
rect 179505 141538 179571 141541
rect 118252 141536 179571 141538
rect 118252 141480 179510 141536
rect 179566 141480 179571 141536
rect 118252 141478 179571 141480
rect 118252 141476 118258 141478
rect 179505 141475 179571 141478
rect 183369 141538 183435 141541
rect 196382 141538 196388 141540
rect 183369 141536 196388 141538
rect 183369 141480 183374 141536
rect 183430 141480 196388 141536
rect 183369 141478 196388 141480
rect 183369 141475 183435 141478
rect 196382 141476 196388 141478
rect 196452 141476 196458 141540
rect 580441 141538 580507 141541
rect 583520 141538 584960 141628
rect 580441 141536 584960 141538
rect 580441 141480 580446 141536
rect 580502 141480 584960 141536
rect 580441 141478 584960 141480
rect 580441 141475 580507 141478
rect 116710 141340 116716 141404
rect 116780 141402 116786 141404
rect 179597 141402 179663 141405
rect 116780 141400 179663 141402
rect 116780 141344 179602 141400
rect 179658 141344 179663 141400
rect 116780 141342 179663 141344
rect 116780 141340 116786 141342
rect 179597 141339 179663 141342
rect 181478 141340 181484 141404
rect 181548 141402 181554 141404
rect 194542 141402 194548 141404
rect 181548 141342 194548 141402
rect 181548 141340 181554 141342
rect 194542 141340 194548 141342
rect 194612 141340 194618 141404
rect 583520 141388 584960 141478
rect -960 140858 480 140948
rect 3509 140858 3575 140861
rect -960 140856 3575 140858
rect -960 140800 3514 140856
rect 3570 140800 3575 140856
rect -960 140798 3575 140800
rect -960 140708 480 140798
rect 3509 140795 3575 140798
rect 120942 140660 120948 140724
rect 121012 140722 121018 140724
rect 137277 140722 137343 140725
rect 121012 140720 137343 140722
rect 121012 140664 137282 140720
rect 137338 140664 137343 140720
rect 121012 140662 137343 140664
rect 121012 140660 121018 140662
rect 137277 140659 137343 140662
rect 184841 140722 184907 140725
rect 197905 140722 197971 140725
rect 184841 140720 197971 140722
rect 184841 140664 184846 140720
rect 184902 140664 197910 140720
rect 197966 140664 197971 140720
rect 184841 140662 197971 140664
rect 184841 140659 184907 140662
rect 197905 140659 197971 140662
rect 115606 140524 115612 140588
rect 115676 140586 115682 140588
rect 132125 140586 132191 140589
rect 115676 140584 132191 140586
rect 115676 140528 132130 140584
rect 132186 140528 132191 140584
rect 115676 140526 132191 140528
rect 115676 140524 115682 140526
rect 132125 140523 132191 140526
rect 183277 140586 183343 140589
rect 193622 140586 193628 140588
rect 183277 140584 193628 140586
rect 183277 140528 183282 140584
rect 183338 140528 193628 140584
rect 183277 140526 193628 140528
rect 183277 140523 183343 140526
rect 193622 140524 193628 140526
rect 193692 140524 193698 140588
rect 113582 140388 113588 140452
rect 113652 140450 113658 140452
rect 130469 140450 130535 140453
rect 113652 140448 130535 140450
rect 113652 140392 130474 140448
rect 130530 140392 130535 140448
rect 113652 140390 130535 140392
rect 113652 140388 113658 140390
rect 130469 140387 130535 140390
rect 186129 140450 186195 140453
rect 192569 140450 192635 140453
rect 186129 140448 192635 140450
rect 186129 140392 186134 140448
rect 186190 140392 192574 140448
rect 192630 140392 192635 140448
rect 186129 140390 192635 140392
rect 186129 140387 186195 140390
rect 192569 140387 192635 140390
rect 115381 140314 115447 140317
rect 134374 140314 134380 140316
rect 115381 140312 134380 140314
rect 115381 140256 115386 140312
rect 115442 140256 134380 140312
rect 115381 140254 134380 140256
rect 115381 140251 115447 140254
rect 134374 140252 134380 140254
rect 134444 140252 134450 140316
rect 179229 140314 179295 140317
rect 194726 140314 194732 140316
rect 179229 140312 194732 140314
rect 179229 140256 179234 140312
rect 179290 140256 194732 140312
rect 179229 140254 194732 140256
rect 179229 140251 179295 140254
rect 194726 140252 194732 140254
rect 194796 140252 194802 140316
rect 120574 140116 120580 140180
rect 120644 140178 120650 140180
rect 141509 140178 141575 140181
rect 120644 140176 141575 140178
rect 120644 140120 141514 140176
rect 141570 140120 141575 140176
rect 120644 140118 141575 140120
rect 120644 140116 120650 140118
rect 141509 140115 141575 140118
rect 162761 140178 162827 140181
rect 187366 140178 187372 140180
rect 162761 140176 187372 140178
rect 162761 140120 162766 140176
rect 162822 140120 187372 140176
rect 162761 140118 187372 140120
rect 162761 140115 162827 140118
rect 187366 140116 187372 140118
rect 187436 140116 187442 140180
rect 121862 139980 121868 140044
rect 121932 140042 121938 140044
rect 147305 140042 147371 140045
rect 121932 140040 147371 140042
rect 121932 139984 147310 140040
rect 147366 139984 147371 140040
rect 121932 139982 147371 139984
rect 121932 139980 121938 139982
rect 147305 139979 147371 139982
rect 154389 140042 154455 140045
rect 188102 140042 188108 140044
rect 154389 140040 188108 140042
rect 154389 139984 154394 140040
rect 154450 139984 188108 140040
rect 154389 139982 188108 139984
rect 154389 139979 154455 139982
rect 188102 139980 188108 139982
rect 188172 139980 188178 140044
rect 188889 140042 188955 140045
rect 196198 140042 196204 140044
rect 188889 140040 196204 140042
rect 188889 139984 188894 140040
rect 188950 139984 196204 140040
rect 188889 139982 196204 139984
rect 188889 139979 188955 139982
rect 196198 139980 196204 139982
rect 196268 139980 196274 140044
rect 115422 139844 115428 139908
rect 115492 139906 115498 139908
rect 124305 139906 124371 139909
rect 115492 139904 124371 139906
rect 115492 139848 124310 139904
rect 124366 139848 124371 139904
rect 115492 139846 124371 139848
rect 115492 139844 115498 139846
rect 124305 139843 124371 139846
rect 187141 139770 187207 139773
rect 187550 139770 187556 139772
rect 187141 139768 187556 139770
rect 187141 139712 187146 139768
rect 187202 139712 187556 139768
rect 187141 139710 187556 139712
rect 187141 139707 187207 139710
rect 187550 139708 187556 139710
rect 187620 139708 187626 139772
rect 125869 139634 125935 139637
rect 187417 139634 187483 139637
rect 122054 139632 125935 139634
rect 122054 139576 125874 139632
rect 125930 139576 125935 139632
rect 122054 139574 125935 139576
rect 116894 139436 116900 139500
rect 116964 139498 116970 139500
rect 117129 139498 117195 139501
rect 122054 139498 122114 139574
rect 125869 139571 125935 139574
rect 187374 139632 187483 139634
rect 187374 139576 187422 139632
rect 187478 139576 187483 139632
rect 187374 139571 187483 139576
rect 124121 139498 124187 139501
rect 116964 139496 117195 139498
rect 116964 139440 117134 139496
rect 117190 139440 117195 139496
rect 116964 139438 117195 139440
rect 116964 139436 116970 139438
rect 117129 139435 117195 139438
rect 121870 139438 122114 139498
rect 123710 139496 124187 139498
rect 123710 139440 124126 139496
rect 124182 139440 124187 139496
rect 123710 139438 124187 139440
rect 121870 139362 121930 139438
rect 118650 139302 121930 139362
rect 108205 139090 108271 139093
rect 118650 139090 118710 139302
rect 122046 139300 122052 139364
rect 122116 139362 122122 139364
rect 123710 139362 123770 139438
rect 124121 139435 124187 139438
rect 182173 139498 182239 139501
rect 186313 139498 186379 139501
rect 182173 139496 182282 139498
rect 182173 139440 182178 139496
rect 182234 139440 182282 139496
rect 182173 139435 182282 139440
rect 122116 139302 123770 139362
rect 122116 139300 122122 139302
rect 123886 139300 123892 139364
rect 123956 139362 123962 139364
rect 124029 139362 124095 139365
rect 125961 139362 126027 139365
rect 123956 139360 124095 139362
rect 123956 139304 124034 139360
rect 124090 139304 124095 139360
rect 123956 139302 124095 139304
rect 123956 139300 123962 139302
rect 124029 139299 124095 139302
rect 124630 139360 126027 139362
rect 124630 139304 125966 139360
rect 126022 139304 126027 139360
rect 124630 139302 126027 139304
rect 108205 139088 118710 139090
rect 108205 139032 108210 139088
rect 108266 139032 118710 139088
rect 108205 139030 118710 139032
rect 120625 139090 120691 139093
rect 124630 139090 124690 139302
rect 125961 139299 126027 139302
rect 126094 139300 126100 139364
rect 126164 139362 126170 139364
rect 128445 139362 128511 139365
rect 126164 139360 128511 139362
rect 126164 139304 128450 139360
rect 128506 139304 128511 139360
rect 126164 139302 128511 139304
rect 126164 139300 126170 139302
rect 128445 139299 128511 139302
rect 136950 139300 136956 139364
rect 137020 139362 137026 139364
rect 141601 139362 141667 139365
rect 146661 139362 146727 139365
rect 154021 139362 154087 139365
rect 137020 139360 141667 139362
rect 137020 139304 141606 139360
rect 141662 139304 141667 139360
rect 137020 139302 141667 139304
rect 137020 139300 137026 139302
rect 141601 139299 141667 139302
rect 142110 139360 146727 139362
rect 142110 139304 146666 139360
rect 146722 139304 146727 139360
rect 142110 139302 146727 139304
rect 120625 139088 124690 139090
rect 120625 139032 120630 139088
rect 120686 139032 124690 139088
rect 120625 139030 124690 139032
rect 108205 139027 108271 139030
rect 120625 139027 120691 139030
rect 115197 138954 115263 138957
rect 142110 138954 142170 139302
rect 146661 139299 146727 139302
rect 151770 139360 154087 139362
rect 151770 139304 154026 139360
rect 154082 139304 154087 139360
rect 151770 139302 154087 139304
rect 115197 138952 142170 138954
rect 115197 138896 115202 138952
rect 115258 138896 142170 138952
rect 115197 138894 142170 138896
rect 115197 138891 115263 138894
rect 108246 138756 108252 138820
rect 108316 138818 108322 138820
rect 136950 138818 136956 138820
rect 108316 138758 136956 138818
rect 108316 138756 108322 138758
rect 136950 138756 136956 138758
rect 137020 138756 137026 138820
rect 119889 138682 119955 138685
rect 151770 138682 151830 139302
rect 154021 139299 154087 139302
rect 180517 139362 180583 139365
rect 180701 139362 180767 139365
rect 180517 139360 180626 139362
rect 180517 139304 180522 139360
rect 180578 139304 180626 139360
rect 180517 139299 180626 139304
rect 180701 139360 182098 139362
rect 180701 139304 180706 139360
rect 180762 139304 182098 139360
rect 180701 139302 182098 139304
rect 180701 139299 180767 139302
rect 180566 138818 180626 139299
rect 182038 138818 182098 139302
rect 182222 138954 182282 139435
rect 186270 139496 186379 139498
rect 186270 139440 186318 139496
rect 186374 139440 186379 139496
rect 186270 139435 186379 139440
rect 186270 139090 186330 139435
rect 186405 139362 186471 139365
rect 187049 139362 187115 139365
rect 187182 139362 187188 139364
rect 186405 139360 186514 139362
rect 186405 139304 186410 139360
rect 186466 139304 186514 139360
rect 186405 139299 186514 139304
rect 187049 139360 187188 139362
rect 187049 139304 187054 139360
rect 187110 139304 187188 139360
rect 187049 139302 187188 139304
rect 187049 139299 187115 139302
rect 187182 139300 187188 139302
rect 187252 139300 187258 139364
rect 186454 139226 186514 139299
rect 186998 139226 187004 139228
rect 186454 139166 187004 139226
rect 186998 139164 187004 139166
rect 187068 139164 187074 139228
rect 187374 139226 187434 139571
rect 187509 139498 187575 139501
rect 187509 139496 187802 139498
rect 187509 139440 187514 139496
rect 187570 139440 187802 139496
rect 187509 139438 187802 139440
rect 187509 139435 187575 139438
rect 187742 139362 187802 139438
rect 192201 139362 192267 139365
rect 187742 139360 192267 139362
rect 187742 139304 192206 139360
rect 192262 139304 192267 139360
rect 187742 139302 192267 139304
rect 192201 139299 192267 139302
rect 195237 139226 195303 139229
rect 187374 139224 195303 139226
rect 187374 139168 195242 139224
rect 195298 139168 195303 139224
rect 187374 139166 195303 139168
rect 195237 139163 195303 139166
rect 197721 139090 197787 139093
rect 186270 139088 197787 139090
rect 186270 139032 197726 139088
rect 197782 139032 197787 139088
rect 186270 139030 197787 139032
rect 197721 139027 197787 139030
rect 190678 138954 190684 138956
rect 182222 138894 190684 138954
rect 190678 138892 190684 138894
rect 190748 138892 190754 138956
rect 193806 138818 193812 138820
rect 180566 138758 180810 138818
rect 182038 138758 193812 138818
rect 119889 138680 151830 138682
rect 119889 138624 119894 138680
rect 119950 138624 151830 138680
rect 119889 138622 151830 138624
rect 180750 138682 180810 138758
rect 193806 138756 193812 138758
rect 193876 138756 193882 138820
rect 199469 138682 199535 138685
rect 180750 138680 199535 138682
rect 180750 138624 199474 138680
rect 199530 138624 199535 138680
rect 180750 138622 199535 138624
rect 119889 138619 119955 138622
rect 199469 138619 199535 138622
rect 120717 138546 120783 138549
rect 126094 138546 126100 138548
rect 120717 138544 126100 138546
rect 120717 138488 120722 138544
rect 120778 138488 126100 138544
rect 120717 138486 126100 138488
rect 120717 138483 120783 138486
rect 126094 138484 126100 138486
rect 126164 138484 126170 138548
rect 185342 138212 185348 138276
rect 185412 138274 185418 138276
rect 186262 138274 186268 138276
rect 185412 138214 186268 138274
rect 185412 138212 185418 138214
rect 186262 138212 186268 138214
rect 186332 138212 186338 138276
rect 115841 138140 115907 138141
rect 115790 138138 115796 138140
rect 115750 138078 115796 138138
rect 115860 138136 115907 138140
rect 115902 138080 115907 138136
rect 115790 138076 115796 138078
rect 115860 138076 115907 138080
rect 115841 138075 115907 138076
rect 118417 138002 118483 138005
rect 122966 138002 122972 138004
rect 118417 138000 122972 138002
rect 118417 137944 118422 138000
rect 118478 137944 122972 138000
rect 118417 137942 122972 137944
rect 118417 137939 118483 137942
rect 122966 137940 122972 137942
rect 123036 137940 123042 138004
rect 111190 137804 111196 137868
rect 111260 137866 111266 137868
rect 124806 137866 124812 137868
rect 111260 137806 124812 137866
rect 111260 137804 111266 137806
rect 124806 137804 124812 137806
rect 124876 137804 124882 137868
rect 185710 137804 185716 137868
rect 185780 137866 185786 137868
rect 193254 137866 193260 137868
rect 185780 137806 193260 137866
rect 185780 137804 185786 137806
rect 193254 137804 193260 137806
rect 193324 137804 193330 137868
rect 187182 137396 187188 137460
rect 187252 137458 187258 137460
rect 195421 137458 195487 137461
rect 187252 137456 195487 137458
rect 187252 137400 195426 137456
rect 195482 137400 195487 137456
rect 187252 137398 195487 137400
rect 187252 137396 187258 137398
rect 195421 137395 195487 137398
rect 580165 137458 580231 137461
rect 583520 137458 584960 137548
rect 580165 137456 584960 137458
rect 580165 137400 580170 137456
rect 580226 137400 584960 137456
rect 580165 137398 584960 137400
rect 580165 137395 580231 137398
rect 187550 137260 187556 137324
rect 187620 137322 187626 137324
rect 200757 137322 200823 137325
rect 187620 137320 200823 137322
rect 187620 137264 200762 137320
rect 200818 137264 200823 137320
rect 583520 137308 584960 137398
rect 187620 137262 200823 137264
rect 187620 137260 187626 137262
rect 200757 137259 200823 137262
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 186814 136580 186820 136644
rect 186884 136642 186890 136644
rect 189901 136642 189967 136645
rect 186884 136640 189967 136642
rect 186884 136584 189906 136640
rect 189962 136584 189967 136640
rect 186884 136582 189967 136584
rect 186884 136580 186890 136582
rect 189901 136579 189967 136582
rect 186262 134404 186268 134468
rect 186332 134466 186338 134468
rect 200849 134466 200915 134469
rect 186332 134464 200915 134466
rect 186332 134408 200854 134464
rect 200910 134408 200915 134464
rect 186332 134406 200915 134408
rect 186332 134404 186338 134406
rect 200849 134403 200915 134406
rect 580717 133378 580783 133381
rect 583520 133378 584960 133468
rect 580717 133376 584960 133378
rect 580717 133320 580722 133376
rect 580778 133320 584960 133376
rect 580717 133318 584960 133320
rect 580717 133315 580783 133318
rect 583520 133228 584960 133318
rect -960 132548 480 132788
rect 122046 132636 122052 132700
rect 122116 132698 122122 132700
rect 122782 132698 122788 132700
rect 122116 132638 122788 132698
rect 122116 132636 122122 132638
rect 122782 132636 122788 132638
rect 122852 132636 122858 132700
rect 122046 132364 122052 132428
rect 122116 132426 122122 132428
rect 122782 132426 122788 132428
rect 122116 132366 122788 132426
rect 122116 132364 122122 132366
rect 122782 132364 122788 132366
rect 122852 132364 122858 132428
rect 580349 129298 580415 129301
rect 583520 129298 584960 129388
rect 580349 129296 584960 129298
rect 580349 129240 580354 129296
rect 580410 129240 584960 129296
rect 580349 129238 584960 129240
rect 580349 129235 580415 129238
rect 583520 129148 584960 129238
rect -960 128468 480 128708
rect 580165 125218 580231 125221
rect 583520 125218 584960 125308
rect 580165 125216 584960 125218
rect 580165 125160 580170 125216
rect 580226 125160 584960 125216
rect 580165 125158 584960 125160
rect 580165 125155 580231 125158
rect 583520 125068 584960 125158
rect -960 124388 480 124628
rect 122046 122980 122052 123044
rect 122116 123042 122122 123044
rect 122782 123042 122788 123044
rect 122116 122982 122788 123042
rect 122116 122980 122122 122982
rect 122782 122980 122788 122982
rect 122852 122980 122858 123044
rect 121729 122770 121795 122773
rect 122782 122770 122788 122772
rect 121729 122768 122788 122770
rect 121729 122712 121734 122768
rect 121790 122712 122788 122768
rect 121729 122710 122788 122712
rect 121729 122707 121795 122710
rect 122782 122708 122788 122710
rect 122852 122708 122858 122772
rect 580625 121138 580691 121141
rect 583520 121138 584960 121228
rect 580625 121136 584960 121138
rect 580625 121080 580630 121136
rect 580686 121080 584960 121136
rect 580625 121078 584960 121080
rect 580625 121075 580691 121078
rect 583520 120988 584960 121078
rect -960 120458 480 120548
rect 3141 120458 3207 120461
rect -960 120456 3207 120458
rect -960 120400 3146 120456
rect 3202 120400 3207 120456
rect -960 120398 3207 120400
rect -960 120308 480 120398
rect 3141 120395 3207 120398
rect -960 117058 480 117148
rect 3233 117058 3299 117061
rect -960 117056 3299 117058
rect -960 117000 3238 117056
rect 3294 117000 3299 117056
rect -960 116998 3299 117000
rect -960 116908 480 116998
rect 3233 116995 3299 116998
rect 580533 117058 580599 117061
rect 583520 117058 584960 117148
rect 580533 117056 584960 117058
rect 580533 117000 580538 117056
rect 580594 117000 584960 117056
rect 580533 116998 584960 117000
rect 580533 116995 580599 116998
rect 583520 116908 584960 116998
rect 121729 113250 121795 113253
rect 122782 113250 122788 113252
rect 121729 113248 122788 113250
rect 121729 113192 121734 113248
rect 121790 113192 122788 113248
rect 121729 113190 122788 113192
rect 121729 113187 121795 113190
rect 122782 113188 122788 113190
rect 122852 113188 122858 113252
rect 121729 113114 121795 113117
rect 122782 113114 122788 113116
rect 121729 113112 122788 113114
rect -960 112978 480 113068
rect 121729 113056 121734 113112
rect 121790 113056 122788 113112
rect 121729 113054 122788 113056
rect 121729 113051 121795 113054
rect 122782 113052 122788 113054
rect 122852 113052 122858 113116
rect 3417 112978 3483 112981
rect -960 112976 3483 112978
rect -960 112920 3422 112976
rect 3478 112920 3483 112976
rect -960 112918 3483 112920
rect -960 112828 480 112918
rect 3417 112915 3483 112918
rect 580165 112978 580231 112981
rect 583520 112978 584960 113068
rect 580165 112976 584960 112978
rect 580165 112920 580170 112976
rect 580226 112920 584960 112976
rect 580165 112918 584960 112920
rect 580165 112915 580231 112918
rect 583520 112828 584960 112918
rect -960 108898 480 108988
rect 3417 108898 3483 108901
rect -960 108896 3483 108898
rect -960 108840 3422 108896
rect 3478 108840 3483 108896
rect -960 108838 3483 108840
rect -960 108748 480 108838
rect 3417 108835 3483 108838
rect 580441 108898 580507 108901
rect 583520 108898 584960 108988
rect 580441 108896 584960 108898
rect 580441 108840 580446 108896
rect 580502 108840 584960 108896
rect 580441 108838 584960 108840
rect 580441 108835 580507 108838
rect 583520 108748 584960 108838
rect -960 104818 480 104908
rect 3417 104818 3483 104821
rect -960 104816 3483 104818
rect -960 104760 3422 104816
rect 3478 104760 3483 104816
rect -960 104758 3483 104760
rect -960 104668 480 104758
rect 3417 104755 3483 104758
rect 580349 104818 580415 104821
rect 583520 104818 584960 104908
rect 580349 104816 584960 104818
rect 580349 104760 580354 104816
rect 580410 104760 584960 104816
rect 580349 104758 584960 104760
rect 580349 104755 580415 104758
rect 583520 104668 584960 104758
rect 121729 103594 121795 103597
rect 122782 103594 122788 103596
rect 121729 103592 122788 103594
rect 121729 103536 121734 103592
rect 121790 103536 122788 103592
rect 121729 103534 122788 103536
rect 121729 103531 121795 103534
rect 122782 103532 122788 103534
rect 122852 103532 122858 103596
rect 121729 103458 121795 103461
rect 122782 103458 122788 103460
rect 121729 103456 122788 103458
rect 121729 103400 121734 103456
rect 121790 103400 122788 103456
rect 121729 103398 122788 103400
rect 121729 103395 121795 103398
rect 122782 103396 122788 103398
rect 122852 103396 122858 103460
rect 580625 101418 580691 101421
rect 583520 101418 584960 101508
rect 580625 101416 584960 101418
rect 580625 101360 580630 101416
rect 580686 101360 584960 101416
rect 580625 101358 584960 101360
rect 580625 101355 580691 101358
rect 583520 101268 584960 101358
rect -960 100738 480 100828
rect 3325 100738 3391 100741
rect -960 100736 3391 100738
rect -960 100680 3330 100736
rect 3386 100680 3391 100736
rect -960 100678 3391 100680
rect -960 100588 480 100678
rect 3325 100675 3391 100678
rect 580441 97338 580507 97341
rect 583520 97338 584960 97428
rect 580441 97336 584960 97338
rect 580441 97280 580446 97336
rect 580502 97280 584960 97336
rect 580441 97278 584960 97280
rect 580441 97275 580507 97278
rect 583520 97188 584960 97278
rect -960 96658 480 96748
rect 3417 96658 3483 96661
rect -960 96656 3483 96658
rect -960 96600 3422 96656
rect 3478 96600 3483 96656
rect -960 96598 3483 96600
rect -960 96508 480 96598
rect 3417 96595 3483 96598
rect 121729 93938 121795 93941
rect 122782 93938 122788 93940
rect 121729 93936 122788 93938
rect 121729 93880 121734 93936
rect 121790 93880 122788 93936
rect 121729 93878 122788 93880
rect 121729 93875 121795 93878
rect 122782 93876 122788 93878
rect 122852 93876 122858 93940
rect 121729 93802 121795 93805
rect 122782 93802 122788 93804
rect 121729 93800 122788 93802
rect 121729 93744 121734 93800
rect 121790 93744 122788 93800
rect 121729 93742 122788 93744
rect 121729 93739 121795 93742
rect 122782 93740 122788 93742
rect 122852 93740 122858 93804
rect 580717 93258 580783 93261
rect 583520 93258 584960 93348
rect 580717 93256 584960 93258
rect 580717 93200 580722 93256
rect 580778 93200 584960 93256
rect 580717 93198 584960 93200
rect 580717 93195 580783 93198
rect 583520 93108 584960 93198
rect -960 92578 480 92668
rect 3141 92578 3207 92581
rect -960 92576 3207 92578
rect -960 92520 3146 92576
rect 3202 92520 3207 92576
rect -960 92518 3207 92520
rect -960 92428 480 92518
rect 3141 92515 3207 92518
rect 115841 92578 115907 92581
rect 120574 92578 120580 92580
rect 115841 92576 120580 92578
rect 115841 92520 115846 92576
rect 115902 92520 120580 92576
rect 115841 92518 120580 92520
rect 115841 92515 115907 92518
rect 120574 92516 120580 92518
rect 120644 92516 120650 92580
rect 186078 91156 186084 91220
rect 186148 91218 186154 91220
rect 188981 91218 189047 91221
rect 186148 91216 189047 91218
rect 186148 91160 188986 91216
rect 189042 91160 189047 91216
rect 186148 91158 189047 91160
rect 186148 91156 186154 91158
rect 188981 91155 189047 91158
rect 580533 89178 580599 89181
rect 583520 89178 584960 89268
rect 580533 89176 584960 89178
rect 580533 89120 580538 89176
rect 580594 89120 584960 89176
rect 580533 89118 584960 89120
rect 580533 89115 580599 89118
rect 583520 89028 584960 89118
rect -960 88348 480 88588
rect 580165 85098 580231 85101
rect 583520 85098 584960 85188
rect 580165 85096 584960 85098
rect 580165 85040 580170 85096
rect 580226 85040 584960 85096
rect 580165 85038 584960 85040
rect 580165 85035 580231 85038
rect 583520 84948 584960 85038
rect -960 84418 480 84508
rect 3417 84418 3483 84421
rect -960 84416 3483 84418
rect -960 84360 3422 84416
rect 3478 84360 3483 84416
rect -960 84358 3483 84360
rect -960 84268 480 84358
rect 3417 84355 3483 84358
rect 111149 83466 111215 83469
rect 122966 83466 122972 83468
rect 111149 83464 122972 83466
rect 111149 83408 111154 83464
rect 111210 83408 122972 83464
rect 111149 83406 122972 83408
rect 111149 83403 111215 83406
rect 122966 83404 122972 83406
rect 123036 83404 123042 83468
rect 187182 82724 187188 82788
rect 187252 82786 187258 82788
rect 191189 82786 191255 82789
rect 187252 82784 191255 82786
rect 187252 82728 191194 82784
rect 191250 82728 191255 82784
rect 187252 82726 191255 82728
rect 187252 82724 187258 82726
rect 191189 82723 191255 82726
rect 186078 82180 186084 82244
rect 186148 82242 186154 82244
rect 193806 82242 193812 82244
rect 186148 82182 193812 82242
rect 186148 82180 186154 82182
rect 193806 82180 193812 82182
rect 193876 82180 193882 82244
rect 100201 81970 100267 81973
rect 135846 81970 135852 81972
rect 100201 81968 135852 81970
rect 100201 81912 100206 81968
rect 100262 81912 135852 81968
rect 100201 81910 135852 81912
rect 100201 81907 100267 81910
rect 135846 81908 135852 81910
rect 135916 81908 135922 81972
rect 176694 81908 176700 81972
rect 176764 81970 176770 81972
rect 216765 81970 216831 81973
rect 176764 81968 216831 81970
rect 176764 81912 216770 81968
rect 216826 81912 216831 81968
rect 176764 81910 216831 81912
rect 176764 81908 176770 81910
rect 216765 81907 216831 81910
rect 102685 81834 102751 81837
rect 137318 81834 137324 81836
rect 102685 81832 137324 81834
rect 102685 81776 102690 81832
rect 102746 81776 137324 81832
rect 102685 81774 137324 81776
rect 102685 81771 102751 81774
rect 137318 81772 137324 81774
rect 137388 81772 137394 81836
rect 175038 81772 175044 81836
rect 175108 81834 175114 81836
rect 200941 81834 201007 81837
rect 175108 81832 201007 81834
rect 175108 81776 200946 81832
rect 201002 81776 201007 81832
rect 175108 81774 201007 81776
rect 175108 81772 175114 81774
rect 200941 81771 201007 81774
rect 111190 81636 111196 81700
rect 111260 81698 111266 81700
rect 111260 81638 125610 81698
rect 111260 81636 111266 81638
rect 115841 81562 115907 81565
rect 119654 81562 119660 81564
rect 115841 81560 119660 81562
rect 115841 81504 115846 81560
rect 115902 81504 119660 81560
rect 115841 81502 119660 81504
rect 115841 81499 115907 81502
rect 119654 81500 119660 81502
rect 119724 81500 119730 81564
rect 125550 81426 125610 81638
rect 184790 81636 184796 81700
rect 184860 81698 184866 81700
rect 205081 81698 205147 81701
rect 184860 81696 205147 81698
rect 184860 81640 205086 81696
rect 205142 81640 205147 81696
rect 184860 81638 205147 81640
rect 184860 81636 184866 81638
rect 205081 81635 205147 81638
rect 141366 81426 141372 81428
rect 125550 81366 141372 81426
rect 141366 81364 141372 81366
rect 141436 81364 141442 81428
rect 189993 81426 190059 81429
rect 196382 81426 196388 81428
rect 189993 81424 196388 81426
rect 189993 81368 189998 81424
rect 190054 81368 196388 81424
rect 189993 81366 196388 81368
rect 189993 81363 190059 81366
rect 196382 81364 196388 81366
rect 196452 81364 196458 81428
rect 108389 81290 108455 81293
rect 131430 81290 131436 81292
rect 108389 81288 131436 81290
rect 108389 81232 108394 81288
rect 108450 81232 131436 81288
rect 108389 81230 131436 81232
rect 108389 81227 108455 81230
rect 131430 81228 131436 81230
rect 131500 81228 131506 81292
rect 166574 81228 166580 81292
rect 166644 81290 166650 81292
rect 199377 81290 199443 81293
rect 207473 81290 207539 81293
rect 166644 81288 199443 81290
rect 166644 81232 199382 81288
rect 199438 81232 199443 81288
rect 166644 81230 199443 81232
rect 166644 81228 166650 81230
rect 199377 81227 199443 81230
rect 200070 81288 207539 81290
rect 200070 81232 207478 81288
rect 207534 81232 207539 81288
rect 200070 81230 207539 81232
rect 99005 81154 99071 81157
rect 133270 81154 133276 81156
rect 99005 81152 133276 81154
rect 99005 81096 99010 81152
rect 99066 81096 133276 81152
rect 99005 81094 133276 81096
rect 99005 81091 99071 81094
rect 133270 81092 133276 81094
rect 133340 81092 133346 81156
rect 174854 81092 174860 81156
rect 174924 81154 174930 81156
rect 200070 81154 200130 81230
rect 207473 81227 207539 81230
rect 174924 81094 200130 81154
rect 202873 81154 202939 81157
rect 203558 81154 203564 81156
rect 202873 81152 203564 81154
rect 202873 81096 202878 81152
rect 202934 81096 203564 81152
rect 202873 81094 203564 81096
rect 174924 81092 174930 81094
rect 202873 81091 202939 81094
rect 203558 81092 203564 81094
rect 203628 81092 203634 81156
rect 101489 81018 101555 81021
rect 135478 81018 135484 81020
rect 101489 81016 135484 81018
rect 101489 80960 101494 81016
rect 101550 80960 135484 81016
rect 101489 80958 135484 80960
rect 101489 80955 101555 80958
rect 135478 80956 135484 80958
rect 135548 80956 135554 81020
rect 166942 80956 166948 81020
rect 167012 81018 167018 81020
rect 203425 81018 203491 81021
rect 167012 81016 203491 81018
rect 167012 80960 203430 81016
rect 203486 80960 203491 81016
rect 167012 80958 203491 80960
rect 167012 80956 167018 80958
rect 203425 80955 203491 80958
rect 112478 80820 112484 80884
rect 112548 80882 112554 80884
rect 147438 80882 147444 80884
rect 112548 80822 147444 80882
rect 112548 80820 112554 80822
rect 147438 80820 147444 80822
rect 147508 80820 147514 80884
rect 154798 80820 154804 80884
rect 154868 80882 154874 80884
rect 193949 80882 194015 80885
rect 154868 80880 194015 80882
rect 154868 80824 193954 80880
rect 194010 80824 194015 80880
rect 583520 80868 584960 81108
rect 154868 80822 194015 80824
rect 154868 80820 154874 80822
rect 193949 80819 194015 80822
rect 99046 80684 99052 80748
rect 99116 80746 99122 80748
rect 134374 80746 134380 80748
rect 99116 80686 134380 80746
rect 99116 80684 99122 80686
rect 134374 80684 134380 80686
rect 134444 80684 134450 80748
rect 217409 80746 217475 80749
rect 153150 80744 217475 80746
rect 153150 80688 217414 80744
rect 217470 80688 217475 80744
rect 153150 80686 217475 80688
rect 116526 80548 116532 80612
rect 116596 80610 116602 80612
rect 123477 80610 123543 80613
rect 116596 80608 123543 80610
rect 116596 80552 123482 80608
rect 123538 80552 123543 80608
rect 116596 80550 123543 80552
rect 116596 80548 116602 80550
rect 123477 80547 123543 80550
rect -960 80338 480 80428
rect 3417 80338 3483 80341
rect -960 80336 3483 80338
rect -960 80280 3422 80336
rect 3478 80280 3483 80336
rect -960 80278 3483 80280
rect -960 80188 480 80278
rect 3417 80275 3483 80278
rect 131849 80338 131915 80341
rect 131849 80336 139778 80338
rect 131849 80280 131854 80336
rect 131910 80280 139778 80336
rect 131849 80278 139778 80280
rect 131849 80275 131915 80278
rect 132217 80202 132283 80205
rect 132217 80200 133890 80202
rect 132217 80144 132222 80200
rect 132278 80144 133890 80200
rect 132217 80142 133890 80144
rect 132217 80139 132283 80142
rect 131430 80004 131436 80068
rect 131500 80066 131506 80068
rect 131849 80066 131915 80069
rect 131500 80064 131915 80066
rect 131500 80008 131854 80064
rect 131910 80008 131915 80064
rect 131500 80006 131915 80008
rect 131500 80004 131506 80006
rect 131849 80003 131915 80006
rect 132631 79962 132697 79967
rect 132631 79906 132636 79962
rect 132692 79906 132697 79962
rect 132631 79901 132697 79906
rect 133183 79964 133249 79967
rect 133183 79962 133292 79964
rect 133183 79906 133188 79962
rect 133244 79932 133292 79962
rect 133244 79906 133276 79932
rect 133183 79901 133276 79906
rect 127433 79794 127499 79797
rect 132634 79794 132694 79901
rect 133232 79870 133276 79901
rect 133270 79868 133276 79870
rect 133340 79868 133346 79932
rect 127433 79792 132694 79794
rect 127433 79736 127438 79792
rect 127494 79736 132694 79792
rect 127433 79734 132694 79736
rect 132815 79792 132881 79797
rect 132815 79736 132820 79792
rect 132876 79736 132881 79792
rect 127433 79731 127499 79734
rect 132815 79731 132881 79736
rect 132818 79661 132878 79731
rect 128997 79658 129063 79661
rect 132493 79658 132559 79661
rect 128997 79656 132559 79658
rect 128997 79600 129002 79656
rect 129058 79600 132498 79656
rect 132554 79600 132559 79656
rect 128997 79598 132559 79600
rect 132818 79656 132927 79661
rect 132818 79600 132866 79656
rect 132922 79600 132927 79656
rect 132818 79598 132927 79600
rect 133830 79658 133890 80142
rect 139718 79967 139778 80278
rect 153150 80202 153210 80686
rect 217409 80683 217475 80686
rect 177246 80548 177252 80612
rect 177316 80610 177322 80612
rect 177941 80610 178007 80613
rect 177316 80608 178007 80610
rect 177316 80552 177946 80608
rect 178002 80552 178007 80608
rect 177316 80550 178007 80552
rect 177316 80548 177322 80550
rect 177941 80547 178007 80550
rect 186313 80610 186379 80613
rect 190678 80610 190684 80612
rect 186313 80608 190684 80610
rect 186313 80552 186318 80608
rect 186374 80552 190684 80608
rect 186313 80550 190684 80552
rect 186313 80547 186379 80550
rect 190678 80548 190684 80550
rect 190748 80548 190754 80612
rect 179229 80474 179295 80477
rect 185577 80474 185643 80477
rect 179229 80472 185643 80474
rect 179229 80416 179234 80472
rect 179290 80416 185582 80472
rect 185638 80416 185643 80472
rect 179229 80414 185643 80416
rect 179229 80411 179295 80414
rect 185577 80411 185643 80414
rect 188429 80474 188495 80477
rect 189993 80474 190059 80477
rect 188429 80472 190059 80474
rect 188429 80416 188434 80472
rect 188490 80416 189998 80472
rect 190054 80416 190059 80472
rect 188429 80414 190059 80416
rect 188429 80411 188495 80414
rect 189993 80411 190059 80414
rect 154246 80202 154252 80204
rect 151356 80142 153210 80202
rect 153886 80142 154252 80202
rect 151356 80066 151416 80142
rect 149792 80006 151416 80066
rect 149792 79967 149852 80006
rect 153886 79967 153946 80142
rect 154246 80140 154252 80142
rect 154316 80140 154322 80204
rect 161054 80202 161060 80204
rect 154438 80142 161060 80202
rect 154438 79967 154498 80142
rect 161054 80140 161060 80142
rect 161124 80140 161130 80204
rect 169150 80202 169156 80204
rect 166030 80142 169156 80202
rect 166030 79967 166090 80142
rect 169150 80140 169156 80142
rect 169220 80140 169226 80204
rect 188613 80202 188679 80205
rect 169296 80200 188679 80202
rect 169296 80144 188618 80200
rect 188674 80144 188679 80200
rect 169296 80142 188679 80144
rect 169296 79967 169356 80142
rect 188613 80139 188679 80142
rect 179597 80066 179663 80069
rect 186814 80066 186820 80068
rect 179597 80064 186820 80066
rect 179597 80008 179602 80064
rect 179658 80008 186820 80064
rect 179597 80006 186820 80008
rect 179597 80003 179663 80006
rect 186814 80004 186820 80006
rect 186884 80004 186890 80068
rect 134655 79964 134721 79967
rect 134655 79962 134856 79964
rect 134011 79928 134077 79933
rect 134379 79932 134445 79933
rect 134374 79930 134380 79932
rect 134011 79872 134016 79928
rect 134072 79872 134077 79928
rect 134011 79867 134077 79872
rect 134288 79870 134380 79930
rect 134374 79868 134380 79870
rect 134444 79868 134450 79932
rect 134655 79906 134660 79962
rect 134716 79906 134856 79962
rect 136403 79962 136469 79967
rect 135115 79932 135181 79933
rect 135110 79930 135116 79932
rect 134655 79904 134856 79906
rect 134655 79901 134721 79904
rect 134379 79867 134445 79868
rect 134014 79794 134074 79867
rect 134333 79794 134399 79797
rect 134014 79792 134399 79794
rect 134014 79736 134338 79792
rect 134394 79736 134399 79792
rect 134014 79734 134399 79736
rect 134333 79731 134399 79734
rect 134655 79794 134721 79797
rect 134796 79794 134856 79904
rect 135024 79870 135116 79930
rect 135110 79868 135116 79870
rect 135180 79868 135186 79932
rect 135662 79868 135668 79932
rect 135732 79930 135738 79932
rect 135851 79930 135917 79933
rect 136403 79932 136408 79962
rect 136464 79932 136469 79962
rect 136679 79964 136745 79967
rect 136679 79962 136880 79964
rect 135732 79928 135917 79930
rect 135732 79872 135856 79928
rect 135912 79872 135917 79928
rect 135732 79870 135917 79872
rect 135732 79868 135738 79870
rect 135115 79867 135181 79868
rect 135851 79867 135917 79870
rect 136398 79868 136404 79932
rect 136468 79930 136474 79932
rect 136468 79870 136526 79930
rect 136679 79906 136684 79962
rect 136740 79906 136880 79962
rect 136679 79904 136880 79906
rect 136679 79901 136745 79904
rect 136468 79868 136474 79870
rect 136587 79826 136653 79831
rect 134931 79796 134997 79797
rect 135299 79796 135365 79797
rect 135897 79796 135963 79797
rect 134655 79792 134856 79794
rect 134655 79736 134660 79792
rect 134716 79736 134856 79792
rect 134655 79734 134856 79736
rect 134655 79731 134721 79734
rect 134926 79732 134932 79796
rect 134996 79794 135002 79796
rect 135294 79794 135300 79796
rect 134996 79734 135088 79794
rect 135208 79734 135300 79794
rect 134996 79732 135002 79734
rect 135294 79732 135300 79734
rect 135364 79732 135370 79796
rect 135846 79732 135852 79796
rect 135916 79794 135963 79796
rect 135916 79792 136008 79794
rect 135958 79736 136008 79792
rect 135916 79734 136008 79736
rect 135916 79732 135963 79734
rect 136214 79732 136220 79796
rect 136284 79794 136290 79796
rect 136587 79794 136592 79826
rect 136284 79770 136592 79794
rect 136648 79770 136653 79826
rect 136284 79765 136653 79770
rect 136284 79734 136650 79765
rect 136284 79732 136290 79734
rect 134931 79731 134997 79732
rect 135299 79731 135365 79732
rect 135897 79731 135963 79732
rect 136820 79658 136880 79904
rect 136955 79962 137021 79967
rect 136955 79906 136960 79962
rect 137016 79906 137021 79962
rect 137323 79964 137389 79967
rect 137323 79962 137446 79964
rect 137323 79932 137328 79962
rect 137384 79932 137446 79962
rect 136955 79901 137021 79906
rect 133830 79598 136880 79658
rect 136958 79658 137018 79901
rect 137318 79868 137324 79932
rect 137388 79904 137446 79932
rect 137507 79962 137573 79967
rect 137507 79906 137512 79962
rect 137568 79906 137573 79962
rect 137388 79868 137394 79904
rect 137507 79901 137573 79906
rect 137691 79962 137757 79967
rect 137691 79906 137696 79962
rect 137752 79906 137757 79962
rect 137691 79901 137757 79906
rect 138243 79962 138309 79967
rect 138243 79906 138248 79962
rect 138304 79906 138309 79962
rect 138243 79901 138309 79906
rect 138427 79962 138493 79967
rect 138427 79906 138432 79962
rect 138488 79906 138493 79962
rect 138611 79962 138677 79967
rect 138611 79932 138616 79962
rect 138672 79932 138677 79962
rect 139715 79962 139781 79967
rect 138427 79901 138493 79906
rect 137185 79658 137251 79661
rect 136958 79656 137251 79658
rect 136958 79600 137190 79656
rect 137246 79600 137251 79656
rect 136958 79598 137251 79600
rect 128997 79595 129063 79598
rect 132493 79595 132559 79598
rect 132861 79595 132927 79598
rect 137185 79595 137251 79598
rect 102961 79522 103027 79525
rect 137510 79522 137570 79901
rect 137694 79797 137754 79901
rect 137967 79894 138033 79899
rect 137967 79838 137972 79894
rect 138028 79838 138033 79894
rect 137967 79833 138033 79838
rect 137645 79792 137754 79797
rect 137645 79736 137650 79792
rect 137706 79736 137754 79792
rect 137645 79734 137754 79736
rect 137645 79731 137711 79734
rect 137737 79658 137803 79661
rect 137970 79658 138030 79833
rect 138246 79797 138306 79901
rect 138246 79792 138355 79797
rect 138246 79736 138294 79792
rect 138350 79736 138355 79792
rect 138246 79734 138355 79736
rect 138289 79731 138355 79734
rect 137737 79656 138030 79658
rect 137737 79600 137742 79656
rect 137798 79600 138030 79656
rect 137737 79598 138030 79600
rect 138430 79661 138490 79901
rect 138606 79868 138612 79932
rect 138676 79930 138682 79932
rect 139255 79930 139321 79933
rect 138676 79870 138734 79930
rect 138798 79928 139321 79930
rect 138798 79872 139260 79928
rect 139316 79872 139321 79928
rect 138798 79870 139321 79872
rect 138676 79868 138682 79870
rect 138430 79656 138539 79661
rect 138430 79600 138478 79656
rect 138534 79600 138539 79656
rect 138430 79598 138539 79600
rect 137737 79595 137803 79598
rect 138473 79595 138539 79598
rect 138657 79658 138723 79661
rect 138798 79658 138858 79870
rect 139255 79867 139321 79870
rect 139439 79930 139505 79933
rect 139439 79928 139640 79930
rect 139439 79872 139444 79928
rect 139500 79872 139640 79928
rect 139715 79906 139720 79962
rect 139776 79906 139781 79962
rect 140267 79962 140333 79967
rect 140083 79932 140149 79933
rect 140267 79932 140272 79962
rect 140328 79932 140333 79962
rect 143487 79962 143553 79967
rect 140078 79930 140084 79932
rect 139715 79901 139781 79906
rect 139439 79870 139640 79872
rect 139992 79870 140084 79930
rect 139439 79867 139505 79870
rect 139163 79792 139229 79797
rect 139163 79736 139168 79792
rect 139224 79736 139229 79792
rect 139163 79731 139229 79736
rect 139301 79796 139367 79797
rect 139301 79792 139348 79796
rect 139412 79794 139418 79796
rect 139301 79736 139306 79792
rect 139301 79732 139348 79736
rect 139412 79734 139458 79794
rect 139412 79732 139418 79734
rect 139301 79731 139367 79732
rect 138657 79656 138858 79658
rect 138657 79600 138662 79656
rect 138718 79600 138858 79656
rect 138657 79598 138858 79600
rect 138657 79595 138723 79598
rect 102961 79520 137570 79522
rect 102961 79464 102966 79520
rect 103022 79464 137570 79520
rect 102961 79462 137570 79464
rect 102961 79459 103027 79462
rect 138054 79460 138060 79524
rect 138124 79522 138130 79524
rect 139166 79522 139226 79731
rect 138124 79462 139226 79522
rect 138124 79460 138130 79462
rect 122414 79324 122420 79388
rect 122484 79386 122490 79388
rect 138381 79386 138447 79389
rect 138606 79386 138612 79388
rect 122484 79326 138030 79386
rect 122484 79324 122490 79326
rect 105813 79250 105879 79253
rect 137369 79250 137435 79253
rect 105813 79248 137435 79250
rect 105813 79192 105818 79248
rect 105874 79192 137374 79248
rect 137430 79192 137435 79248
rect 105813 79190 137435 79192
rect 105813 79187 105879 79190
rect 137369 79187 137435 79190
rect 101581 79114 101647 79117
rect 135110 79114 135116 79116
rect 101581 79112 135116 79114
rect 101581 79056 101586 79112
rect 101642 79056 135116 79112
rect 101581 79054 135116 79056
rect 101581 79051 101647 79054
rect 135110 79052 135116 79054
rect 135180 79052 135186 79116
rect 135478 79052 135484 79116
rect 135548 79114 135554 79116
rect 135621 79114 135687 79117
rect 135548 79112 135687 79114
rect 135548 79056 135626 79112
rect 135682 79056 135687 79112
rect 135548 79054 135687 79056
rect 135548 79052 135554 79054
rect 135621 79051 135687 79054
rect 136633 79114 136699 79117
rect 136766 79114 136772 79116
rect 136633 79112 136772 79114
rect 136633 79056 136638 79112
rect 136694 79056 136772 79112
rect 136633 79054 136772 79056
rect 136633 79051 136699 79054
rect 136766 79052 136772 79054
rect 136836 79052 136842 79116
rect 102869 78978 102935 78981
rect 137461 78978 137527 78981
rect 102869 78976 137527 78978
rect 102869 78920 102874 78976
rect 102930 78920 137466 78976
rect 137522 78920 137527 78976
rect 102869 78918 137527 78920
rect 137970 78978 138030 79326
rect 138381 79384 138612 79386
rect 138381 79328 138386 79384
rect 138442 79328 138612 79384
rect 138381 79326 138612 79328
rect 138381 79323 138447 79326
rect 138606 79324 138612 79326
rect 138676 79324 138682 79388
rect 139117 79386 139183 79389
rect 139580 79386 139640 79870
rect 140078 79868 140084 79870
rect 140148 79868 140154 79932
rect 140262 79868 140268 79932
rect 140332 79930 140338 79932
rect 140635 79930 140701 79933
rect 140332 79870 140390 79930
rect 140454 79928 140701 79930
rect 140454 79872 140640 79928
rect 140696 79872 140701 79928
rect 140454 79870 140701 79872
rect 140332 79868 140338 79870
rect 140083 79867 140149 79868
rect 139945 79794 140011 79797
rect 140454 79794 140514 79870
rect 140635 79867 140701 79870
rect 140911 79930 140977 79933
rect 141182 79930 141188 79932
rect 140911 79928 141188 79930
rect 140911 79872 140916 79928
rect 140972 79872 141188 79928
rect 140911 79870 141188 79872
rect 140911 79867 140977 79870
rect 141182 79868 141188 79870
rect 141252 79868 141258 79932
rect 142935 79930 143001 79933
rect 141742 79928 143001 79930
rect 141742 79872 142940 79928
rect 142996 79872 143001 79928
rect 143487 79906 143492 79962
rect 143548 79906 143553 79962
rect 145235 79962 145301 79967
rect 143487 79901 143553 79906
rect 141742 79870 143001 79872
rect 139945 79792 140514 79794
rect 139945 79736 139950 79792
rect 140006 79736 140514 79792
rect 139945 79734 140514 79736
rect 139945 79731 140011 79734
rect 140630 79732 140636 79796
rect 140700 79794 140706 79796
rect 141742 79794 141802 79870
rect 142935 79867 143001 79870
rect 143490 79797 143550 79901
rect 144494 79868 144500 79932
rect 144564 79930 144570 79932
rect 144775 79930 144841 79933
rect 144564 79928 144841 79930
rect 144564 79872 144780 79928
rect 144836 79872 144841 79928
rect 145235 79906 145240 79962
rect 145296 79906 145301 79962
rect 145235 79901 145301 79906
rect 145603 79962 145669 79967
rect 145603 79906 145608 79962
rect 145664 79906 145669 79962
rect 145603 79901 145669 79906
rect 145879 79964 145945 79967
rect 145879 79962 145988 79964
rect 145879 79906 145884 79962
rect 145940 79906 145988 79962
rect 145879 79901 145988 79906
rect 146155 79962 146221 79967
rect 146155 79906 146160 79962
rect 146216 79906 146221 79962
rect 147443 79964 147509 79967
rect 147443 79962 147566 79964
rect 147075 79930 147141 79933
rect 147443 79932 147448 79962
rect 147504 79932 147566 79962
rect 146155 79901 146221 79906
rect 146756 79928 147141 79930
rect 144564 79870 144841 79872
rect 144564 79868 144570 79870
rect 144775 79867 144841 79870
rect 140700 79734 141802 79794
rect 143487 79792 143553 79797
rect 143487 79736 143492 79792
rect 143548 79736 143553 79792
rect 140700 79732 140706 79734
rect 143487 79731 143553 79736
rect 143717 79794 143783 79797
rect 144269 79794 144335 79797
rect 143717 79792 144335 79794
rect 143717 79736 143722 79792
rect 143778 79736 144274 79792
rect 144330 79736 144335 79792
rect 143717 79734 144335 79736
rect 143717 79731 143783 79734
rect 144269 79731 144335 79734
rect 145238 79661 145298 79901
rect 145606 79661 145666 79901
rect 141417 79660 141483 79661
rect 141366 79596 141372 79660
rect 141436 79658 141483 79660
rect 141436 79656 141528 79658
rect 141478 79600 141528 79656
rect 141436 79598 141528 79600
rect 141436 79596 141483 79598
rect 143942 79596 143948 79660
rect 144012 79658 144018 79660
rect 144821 79658 144887 79661
rect 145097 79660 145163 79661
rect 145046 79658 145052 79660
rect 144012 79656 144887 79658
rect 144012 79600 144826 79656
rect 144882 79600 144887 79656
rect 144012 79598 144887 79600
rect 145006 79598 145052 79658
rect 145116 79656 145163 79660
rect 145158 79600 145163 79656
rect 144012 79596 144018 79598
rect 141417 79595 141483 79596
rect 144821 79595 144887 79598
rect 145046 79596 145052 79598
rect 145116 79596 145163 79600
rect 145238 79656 145347 79661
rect 145238 79600 145286 79656
rect 145342 79600 145347 79656
rect 145238 79598 145347 79600
rect 145097 79595 145163 79596
rect 145281 79595 145347 79598
rect 145557 79656 145666 79661
rect 145557 79600 145562 79656
rect 145618 79600 145666 79656
rect 145557 79598 145666 79600
rect 145557 79595 145623 79598
rect 140773 79522 140839 79525
rect 141233 79522 141299 79525
rect 140773 79520 141299 79522
rect 140773 79464 140778 79520
rect 140834 79464 141238 79520
rect 141294 79464 141299 79520
rect 140773 79462 141299 79464
rect 140773 79459 140839 79462
rect 141233 79459 141299 79462
rect 144821 79522 144887 79525
rect 145928 79522 145988 79901
rect 144821 79520 145988 79522
rect 144821 79464 144826 79520
rect 144882 79464 145988 79520
rect 144821 79462 145988 79464
rect 144821 79459 144887 79462
rect 139117 79384 139640 79386
rect 139117 79328 139122 79384
rect 139178 79328 139640 79384
rect 139117 79326 139640 79328
rect 140129 79386 140195 79389
rect 140681 79386 140747 79389
rect 140129 79384 140747 79386
rect 140129 79328 140134 79384
rect 140190 79328 140686 79384
rect 140742 79328 140747 79384
rect 140129 79326 140747 79328
rect 139117 79323 139183 79326
rect 140129 79323 140195 79326
rect 140681 79323 140747 79326
rect 145465 79386 145531 79389
rect 146158 79386 146218 79901
rect 146339 79894 146405 79899
rect 146339 79838 146344 79894
rect 146400 79838 146405 79894
rect 146339 79833 146405 79838
rect 146756 79872 147080 79928
rect 147136 79872 147141 79928
rect 146756 79870 147141 79872
rect 146342 79661 146402 79833
rect 146293 79656 146402 79661
rect 146293 79600 146298 79656
rect 146354 79600 146402 79656
rect 146293 79598 146402 79600
rect 146293 79595 146359 79598
rect 146756 79525 146816 79870
rect 147075 79867 147141 79870
rect 147438 79868 147444 79932
rect 147508 79904 147566 79932
rect 147627 79962 147693 79967
rect 147627 79906 147632 79962
rect 147688 79906 147693 79962
rect 149467 79962 149533 79967
rect 148547 79932 148613 79933
rect 148542 79930 148548 79932
rect 147508 79868 147514 79904
rect 147627 79901 147693 79906
rect 147630 79797 147690 79901
rect 148456 79870 148548 79930
rect 148542 79868 148548 79870
rect 148612 79868 148618 79932
rect 149099 79930 149165 79933
rect 149467 79932 149472 79962
rect 149528 79932 149533 79962
rect 149743 79962 149852 79967
rect 149099 79928 149208 79930
rect 149099 79872 149104 79928
rect 149160 79872 149208 79928
rect 148547 79867 148613 79868
rect 149099 79867 149208 79872
rect 149462 79868 149468 79932
rect 149532 79930 149538 79932
rect 149532 79870 149590 79930
rect 149743 79906 149748 79962
rect 149804 79906 149852 79962
rect 151491 79962 151557 79967
rect 149743 79904 149852 79906
rect 150019 79928 150085 79933
rect 149743 79901 149809 79904
rect 150019 79872 150024 79928
rect 150080 79872 150085 79928
rect 150663 79930 150729 79933
rect 150934 79930 150940 79932
rect 150663 79928 150940 79930
rect 149532 79868 149538 79870
rect 150019 79867 150085 79872
rect 150203 79894 150269 79899
rect 147581 79792 147690 79797
rect 148271 79826 148337 79831
rect 148271 79794 148276 79826
rect 147581 79736 147586 79792
rect 147642 79736 147690 79792
rect 147581 79734 147690 79736
rect 148044 79770 148276 79794
rect 148332 79770 148337 79826
rect 148044 79765 148337 79770
rect 148044 79734 148334 79765
rect 147581 79731 147647 79734
rect 148044 79661 148104 79734
rect 149148 79661 149208 79867
rect 150022 79797 150082 79867
rect 150203 79838 150208 79894
rect 150264 79838 150269 79894
rect 150203 79833 150269 79838
rect 150387 79894 150453 79899
rect 150387 79838 150392 79894
rect 150448 79838 150453 79894
rect 150663 79872 150668 79928
rect 150724 79872 150940 79928
rect 150663 79870 150940 79872
rect 150663 79867 150729 79870
rect 150934 79868 150940 79870
rect 151004 79868 151010 79932
rect 151215 79930 151281 79933
rect 151172 79928 151281 79930
rect 151172 79872 151220 79928
rect 151276 79872 151281 79928
rect 151491 79906 151496 79962
rect 151552 79906 151557 79962
rect 151491 79901 151557 79906
rect 151859 79962 151925 79967
rect 152135 79964 152201 79967
rect 151859 79906 151864 79962
rect 151920 79906 151925 79962
rect 151859 79901 151925 79906
rect 152092 79962 152201 79964
rect 152092 79906 152140 79962
rect 152196 79906 152201 79962
rect 152092 79901 152201 79906
rect 152319 79964 152385 79967
rect 152319 79962 152428 79964
rect 152319 79906 152324 79962
rect 152380 79906 152428 79962
rect 153331 79962 153397 79967
rect 152595 79932 152661 79933
rect 152590 79930 152596 79932
rect 152319 79901 152428 79906
rect 151172 79867 151281 79872
rect 150387 79833 150453 79838
rect 149973 79792 150082 79797
rect 149973 79736 149978 79792
rect 150034 79736 150082 79792
rect 149973 79734 150082 79736
rect 149973 79731 150039 79734
rect 148041 79656 148107 79661
rect 148041 79600 148046 79656
rect 148102 79600 148107 79656
rect 148041 79595 148107 79600
rect 148225 79658 148291 79661
rect 148961 79658 149027 79661
rect 148225 79656 148472 79658
rect 148225 79600 148230 79656
rect 148286 79600 148472 79656
rect 148225 79598 148472 79600
rect 148225 79595 148291 79598
rect 148412 79525 148472 79598
rect 148550 79656 149027 79658
rect 148550 79600 148966 79656
rect 149022 79600 149027 79656
rect 148550 79598 149027 79600
rect 146753 79520 146819 79525
rect 146753 79464 146758 79520
rect 146814 79464 146819 79520
rect 146753 79459 146819 79464
rect 148409 79520 148475 79525
rect 148409 79464 148414 79520
rect 148470 79464 148475 79520
rect 148409 79459 148475 79464
rect 145465 79384 146218 79386
rect 145465 79328 145470 79384
rect 145526 79328 146218 79384
rect 145465 79326 146218 79328
rect 145465 79323 145531 79326
rect 147806 79324 147812 79388
rect 147876 79386 147882 79388
rect 148550 79386 148610 79598
rect 148961 79595 149027 79598
rect 149145 79656 149211 79661
rect 149145 79600 149150 79656
rect 149206 79600 149211 79656
rect 149145 79595 149211 79600
rect 147876 79326 148610 79386
rect 149513 79386 149579 79389
rect 150206 79386 150266 79833
rect 150390 79661 150450 79833
rect 151172 79796 151232 79867
rect 151118 79732 151124 79796
rect 151188 79734 151232 79796
rect 151188 79732 151194 79734
rect 150341 79656 150450 79661
rect 150341 79600 150346 79656
rect 150402 79600 150450 79656
rect 150341 79598 150450 79600
rect 150341 79595 150407 79598
rect 151353 79522 151419 79525
rect 151494 79522 151554 79901
rect 151862 79661 151922 79901
rect 151629 79656 151695 79661
rect 151629 79600 151634 79656
rect 151690 79600 151695 79656
rect 151629 79595 151695 79600
rect 151862 79656 151971 79661
rect 151862 79600 151910 79656
rect 151966 79600 151971 79656
rect 151862 79598 151971 79600
rect 152092 79658 152152 79901
rect 152368 79797 152428 79901
rect 152504 79870 152596 79930
rect 152590 79868 152596 79870
rect 152660 79868 152666 79932
rect 152774 79868 152780 79932
rect 152844 79930 152850 79932
rect 153055 79930 153121 79933
rect 152844 79928 153121 79930
rect 152844 79872 153060 79928
rect 153116 79872 153121 79928
rect 153331 79906 153336 79962
rect 153392 79906 153397 79962
rect 153331 79901 153397 79906
rect 153515 79962 153581 79967
rect 153515 79906 153520 79962
rect 153576 79906 153581 79962
rect 153699 79962 153765 79967
rect 153699 79932 153704 79962
rect 153760 79932 153765 79962
rect 153883 79962 153949 79967
rect 153515 79901 153581 79906
rect 152844 79870 153121 79872
rect 152844 79868 152850 79870
rect 152595 79867 152661 79868
rect 153055 79867 153121 79870
rect 152365 79792 152431 79797
rect 152365 79736 152370 79792
rect 152426 79736 152431 79792
rect 152365 79731 152431 79736
rect 152503 79794 152569 79797
rect 152503 79792 152612 79794
rect 152503 79736 152508 79792
rect 152564 79736 152612 79792
rect 152503 79731 152612 79736
rect 152552 79661 152612 79731
rect 152273 79658 152339 79661
rect 152092 79656 152339 79658
rect 152092 79600 152278 79656
rect 152334 79600 152339 79656
rect 152092 79598 152339 79600
rect 151905 79595 151971 79598
rect 152273 79595 152339 79598
rect 152549 79656 152615 79661
rect 152549 79600 152554 79656
rect 152610 79600 152615 79656
rect 152549 79595 152615 79600
rect 153334 79658 153394 79901
rect 153518 79794 153578 79901
rect 153694 79868 153700 79932
rect 153764 79930 153770 79932
rect 153764 79870 153822 79930
rect 153883 79906 153888 79962
rect 153944 79906 153949 79962
rect 154435 79962 154501 79967
rect 154711 79964 154777 79967
rect 154067 79932 154133 79933
rect 153883 79901 153949 79906
rect 153764 79868 153770 79870
rect 154062 79868 154068 79932
rect 154132 79930 154138 79932
rect 154132 79870 154224 79930
rect 154435 79906 154440 79962
rect 154496 79906 154501 79962
rect 154435 79901 154501 79906
rect 154668 79962 154777 79964
rect 154668 79906 154716 79962
rect 154772 79906 154777 79962
rect 154668 79901 154777 79906
rect 155171 79962 155237 79967
rect 155171 79906 155176 79962
rect 155232 79906 155237 79962
rect 155171 79901 155237 79906
rect 155539 79962 155605 79967
rect 157839 79964 157905 79967
rect 155539 79906 155544 79962
rect 155600 79906 155605 79962
rect 157704 79962 157905 79964
rect 155539 79901 155605 79906
rect 157563 79928 157629 79933
rect 154132 79868 154138 79870
rect 154067 79867 154133 79868
rect 154246 79794 154252 79796
rect 153518 79734 154252 79794
rect 154246 79732 154252 79734
rect 154316 79732 154322 79796
rect 154668 79794 154728 79901
rect 154530 79734 154728 79794
rect 154021 79658 154087 79661
rect 153334 79656 154087 79658
rect 153334 79600 154026 79656
rect 154082 79600 154087 79656
rect 153334 79598 154087 79600
rect 154021 79595 154087 79598
rect 151353 79520 151554 79522
rect 151353 79464 151358 79520
rect 151414 79464 151554 79520
rect 151353 79462 151554 79464
rect 151353 79459 151419 79462
rect 149513 79384 150266 79386
rect 149513 79328 149518 79384
rect 149574 79328 150266 79384
rect 149513 79326 150266 79328
rect 147876 79324 147882 79326
rect 149513 79323 149579 79326
rect 139301 79252 139367 79253
rect 139301 79250 139348 79252
rect 139256 79248 139348 79250
rect 139256 79192 139306 79248
rect 139256 79190 139348 79192
rect 139301 79188 139348 79190
rect 139412 79188 139418 79252
rect 140773 79250 140839 79253
rect 141233 79250 141299 79253
rect 140773 79248 141299 79250
rect 140773 79192 140778 79248
rect 140834 79192 141238 79248
rect 141294 79192 141299 79248
rect 140773 79190 141299 79192
rect 151632 79250 151692 79595
rect 154530 79522 154590 79734
rect 154757 79660 154823 79661
rect 154757 79658 154804 79660
rect 154712 79656 154804 79658
rect 154712 79600 154762 79656
rect 154712 79598 154804 79600
rect 154757 79596 154804 79598
rect 154868 79596 154874 79660
rect 154757 79595 154823 79596
rect 154757 79522 154823 79525
rect 154530 79520 154823 79522
rect 154530 79464 154762 79520
rect 154818 79464 154823 79520
rect 154530 79462 154823 79464
rect 155174 79522 155234 79901
rect 155542 79658 155602 79901
rect 157563 79872 157568 79928
rect 157624 79872 157629 79928
rect 157563 79867 157629 79872
rect 157704 79906 157844 79962
rect 157900 79906 157905 79962
rect 157704 79904 157905 79906
rect 157149 79658 157215 79661
rect 155542 79656 157215 79658
rect 155542 79600 157154 79656
rect 157210 79600 157215 79656
rect 155542 79598 157215 79600
rect 157566 79658 157626 79867
rect 157704 79794 157764 79904
rect 157839 79901 157905 79904
rect 158207 79962 158273 79967
rect 158207 79906 158212 79962
rect 158268 79930 158273 79962
rect 162071 79962 162137 79967
rect 158268 79906 160432 79930
rect 158207 79901 160432 79906
rect 158210 79870 160432 79901
rect 157885 79794 157951 79797
rect 157704 79792 157951 79794
rect 157704 79736 157890 79792
rect 157946 79736 157951 79792
rect 157704 79734 157951 79736
rect 157885 79731 157951 79734
rect 158161 79794 158227 79797
rect 158851 79796 158917 79797
rect 158478 79794 158484 79796
rect 158161 79792 158484 79794
rect 158161 79736 158166 79792
rect 158222 79736 158484 79792
rect 158161 79734 158484 79736
rect 158161 79731 158227 79734
rect 158478 79732 158484 79734
rect 158548 79732 158554 79796
rect 158846 79794 158852 79796
rect 158760 79734 158852 79794
rect 158846 79732 158852 79734
rect 158916 79732 158922 79796
rect 159265 79794 159331 79797
rect 159582 79794 159588 79796
rect 159265 79792 159588 79794
rect 159265 79736 159270 79792
rect 159326 79736 159588 79792
rect 159265 79734 159588 79736
rect 158851 79731 158917 79732
rect 159265 79731 159331 79734
rect 159582 79732 159588 79734
rect 159652 79732 159658 79796
rect 159265 79658 159331 79661
rect 157566 79656 159331 79658
rect 157566 79600 159270 79656
rect 159326 79600 159331 79656
rect 157566 79598 159331 79600
rect 160372 79658 160432 79870
rect 160502 79868 160508 79932
rect 160572 79930 160578 79932
rect 160967 79930 161033 79933
rect 160572 79928 161033 79930
rect 160572 79872 160972 79928
rect 161028 79872 161033 79928
rect 160572 79870 161033 79872
rect 160572 79868 160578 79870
rect 160967 79867 161033 79870
rect 161151 79930 161217 79933
rect 161790 79930 161796 79932
rect 161151 79928 161796 79930
rect 161151 79872 161156 79928
rect 161212 79872 161796 79928
rect 161151 79870 161796 79872
rect 161151 79867 161217 79870
rect 161790 79868 161796 79870
rect 161860 79868 161866 79932
rect 162071 79906 162076 79962
rect 162132 79930 162137 79962
rect 162899 79962 162965 79967
rect 162342 79930 162348 79932
rect 162132 79906 162348 79930
rect 162071 79901 162348 79906
rect 162074 79870 162348 79901
rect 162342 79868 162348 79870
rect 162412 79868 162418 79932
rect 162899 79906 162904 79962
rect 162960 79906 162965 79962
rect 163451 79962 163517 79967
rect 163451 79932 163456 79962
rect 163512 79932 163517 79962
rect 165107 79962 165173 79967
rect 162899 79901 162965 79906
rect 161519 79794 161585 79797
rect 161933 79794 161999 79797
rect 161519 79792 161999 79794
rect 161519 79736 161524 79792
rect 161580 79736 161938 79792
rect 161994 79736 161999 79792
rect 161519 79734 161999 79736
rect 161519 79731 161585 79734
rect 161933 79731 161999 79734
rect 162902 79661 162962 79901
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 163911 79930 163977 79933
rect 164279 79930 164345 79933
rect 163516 79870 163574 79930
rect 163868 79928 163977 79930
rect 163868 79872 163916 79928
rect 163972 79872 163977 79928
rect 163516 79868 163522 79870
rect 163868 79867 163977 79872
rect 164144 79928 164345 79930
rect 164144 79872 164284 79928
rect 164340 79872 164345 79928
rect 164144 79870 164345 79872
rect 163630 79732 163636 79796
rect 163700 79794 163706 79796
rect 163868 79794 163928 79867
rect 163700 79734 163928 79794
rect 163700 79732 163706 79734
rect 164144 79661 164204 79870
rect 164279 79867 164345 79870
rect 164463 79930 164529 79933
rect 164463 79928 164664 79930
rect 164463 79872 164468 79928
rect 164524 79872 164664 79928
rect 165107 79906 165112 79962
rect 165168 79906 165173 79962
rect 165107 79901 165173 79906
rect 165291 79962 165357 79967
rect 165291 79906 165296 79962
rect 165352 79906 165357 79962
rect 165843 79962 165909 79967
rect 165291 79901 165357 79906
rect 165475 79930 165541 79933
rect 165475 79928 165768 79930
rect 164463 79870 164664 79872
rect 164463 79867 164529 79870
rect 164604 79796 164664 79870
rect 164550 79732 164556 79796
rect 164620 79734 164664 79796
rect 164620 79732 164626 79734
rect 165110 79661 165170 79901
rect 165294 79797 165354 79901
rect 165475 79872 165480 79928
rect 165536 79872 165768 79928
rect 165843 79906 165848 79962
rect 165904 79906 165909 79962
rect 165843 79901 165909 79906
rect 166027 79962 166093 79967
rect 166027 79906 166032 79962
rect 166088 79906 166093 79962
rect 166027 79901 166093 79906
rect 166579 79962 166645 79967
rect 166579 79906 166584 79962
rect 166640 79930 166645 79962
rect 167039 79964 167105 79967
rect 167039 79962 167148 79964
rect 166758 79930 166764 79932
rect 166640 79906 166764 79930
rect 166579 79901 166764 79906
rect 165475 79870 165768 79872
rect 165475 79867 165541 79870
rect 165708 79797 165768 79870
rect 165245 79792 165354 79797
rect 165245 79736 165250 79792
rect 165306 79736 165354 79792
rect 165245 79734 165354 79736
rect 165705 79792 165771 79797
rect 165705 79736 165710 79792
rect 165766 79736 165771 79792
rect 165245 79731 165311 79734
rect 165705 79731 165771 79736
rect 165846 79794 165906 79901
rect 166582 79870 166764 79901
rect 166758 79868 166764 79870
rect 166828 79868 166834 79932
rect 167039 79906 167044 79962
rect 167100 79932 167148 79962
rect 168603 79962 168669 79967
rect 167100 79906 167132 79932
rect 167039 79901 167132 79906
rect 167088 79870 167132 79901
rect 167126 79868 167132 79870
rect 167196 79868 167202 79932
rect 167407 79930 167473 79933
rect 167867 79932 167933 79933
rect 168235 79932 168301 79933
rect 167862 79930 167868 79932
rect 167407 79928 167516 79930
rect 167407 79872 167412 79928
rect 167468 79872 167516 79928
rect 167407 79867 167516 79872
rect 167776 79870 167868 79930
rect 167862 79868 167868 79870
rect 167932 79868 167938 79932
rect 168230 79930 168236 79932
rect 168144 79870 168236 79930
rect 168230 79868 168236 79870
rect 168300 79868 168306 79932
rect 168603 79906 168608 79962
rect 168664 79906 168669 79962
rect 168603 79901 168669 79906
rect 169247 79962 169356 79967
rect 169247 79906 169252 79962
rect 169308 79906 169356 79962
rect 169983 79964 170049 79967
rect 169983 79962 170092 79964
rect 169247 79904 169356 79906
rect 169615 79930 169681 79933
rect 169615 79928 169724 79930
rect 169247 79901 169313 79904
rect 167867 79867 167933 79868
rect 168235 79867 168301 79868
rect 165981 79794 166047 79797
rect 166947 79796 167013 79797
rect 165846 79792 166047 79794
rect 165846 79736 165986 79792
rect 166042 79736 166047 79792
rect 165846 79734 166047 79736
rect 165981 79731 166047 79734
rect 166942 79732 166948 79796
rect 167012 79794 167018 79796
rect 167012 79734 167104 79794
rect 167012 79732 167018 79734
rect 166947 79731 167013 79732
rect 161473 79658 161539 79661
rect 160372 79656 161539 79658
rect 160372 79600 161478 79656
rect 161534 79600 161539 79656
rect 160372 79598 161539 79600
rect 162902 79656 163011 79661
rect 162902 79600 162950 79656
rect 163006 79600 163011 79656
rect 162902 79598 163011 79600
rect 157149 79595 157215 79598
rect 159265 79595 159331 79598
rect 161473 79595 161539 79598
rect 162945 79595 163011 79598
rect 164141 79656 164207 79661
rect 164141 79600 164146 79656
rect 164202 79600 164207 79656
rect 164141 79595 164207 79600
rect 165061 79656 165170 79661
rect 165061 79600 165066 79656
rect 165122 79600 165170 79656
rect 165061 79598 165170 79600
rect 165613 79658 165679 79661
rect 166533 79660 166599 79661
rect 166390 79658 166396 79660
rect 165613 79656 166396 79658
rect 165613 79600 165618 79656
rect 165674 79600 166396 79656
rect 165613 79598 166396 79600
rect 165061 79595 165127 79598
rect 165613 79595 165679 79598
rect 166390 79596 166396 79598
rect 166460 79596 166466 79660
rect 166533 79656 166580 79660
rect 166644 79658 166650 79660
rect 167456 79658 167516 79867
rect 167678 79732 167684 79796
rect 167748 79794 167754 79796
rect 168051 79794 168117 79797
rect 167748 79792 168117 79794
rect 167748 79736 168056 79792
rect 168112 79736 168117 79792
rect 167748 79734 168117 79736
rect 167748 79732 167754 79734
rect 168051 79731 168117 79734
rect 168046 79658 168052 79660
rect 166533 79600 166538 79656
rect 166533 79596 166580 79600
rect 166644 79598 166690 79658
rect 167456 79598 168052 79658
rect 166644 79596 166650 79598
rect 168046 79596 168052 79598
rect 168116 79596 168122 79660
rect 168606 79658 168666 79901
rect 169615 79872 169620 79928
rect 169676 79872 169724 79928
rect 169983 79906 169988 79962
rect 170044 79932 170092 79962
rect 170259 79962 170325 79967
rect 170044 79906 170076 79932
rect 169983 79901 170076 79906
rect 169615 79867 169724 79872
rect 170032 79870 170076 79901
rect 170070 79868 170076 79870
rect 170140 79868 170146 79932
rect 170259 79906 170264 79962
rect 170320 79906 170325 79962
rect 172283 79962 172349 79967
rect 170259 79901 170325 79906
rect 170719 79930 170785 79933
rect 171087 79930 171153 79933
rect 172283 79932 172288 79962
rect 172344 79932 172349 79962
rect 172467 79962 172533 79967
rect 173111 79964 173177 79967
rect 170719 79928 170828 79930
rect 168741 79658 168807 79661
rect 168606 79656 168807 79658
rect 168606 79600 168746 79656
rect 168802 79600 168807 79656
rect 168606 79598 168807 79600
rect 169664 79658 169724 79867
rect 170262 79794 170322 79901
rect 170719 79872 170724 79928
rect 170780 79872 170828 79928
rect 170719 79867 170828 79872
rect 171087 79928 171196 79930
rect 171087 79872 171092 79928
rect 171148 79872 171196 79928
rect 171087 79867 171196 79872
rect 170768 79796 170828 79867
rect 171136 79797 171196 79867
rect 171915 79894 171981 79899
rect 171915 79838 171920 79894
rect 171976 79838 171981 79894
rect 172278 79868 172284 79932
rect 172348 79930 172354 79932
rect 172348 79870 172406 79930
rect 172467 79906 172472 79962
rect 172528 79906 172533 79962
rect 173068 79962 173177 79964
rect 172467 79901 172533 79906
rect 172651 79928 172717 79933
rect 173068 79932 173116 79962
rect 172348 79868 172354 79870
rect 171915 79833 171981 79838
rect 170622 79794 170628 79796
rect 170262 79734 170628 79794
rect 170622 79732 170628 79734
rect 170692 79732 170698 79796
rect 170768 79734 170812 79796
rect 170806 79732 170812 79734
rect 170876 79732 170882 79796
rect 171133 79792 171199 79797
rect 171593 79796 171659 79797
rect 171542 79794 171548 79796
rect 171133 79736 171138 79792
rect 171194 79736 171199 79792
rect 171133 79731 171199 79736
rect 171502 79734 171548 79794
rect 171612 79792 171659 79796
rect 171654 79736 171659 79792
rect 171542 79732 171548 79734
rect 171612 79732 171659 79736
rect 171593 79731 171659 79732
rect 171225 79658 171291 79661
rect 169664 79656 171291 79658
rect 169664 79600 171230 79656
rect 171286 79600 171291 79656
rect 169664 79598 171291 79600
rect 171918 79658 171978 79833
rect 172470 79797 172530 79901
rect 172651 79872 172656 79928
rect 172712 79872 172717 79928
rect 172651 79867 172717 79872
rect 173014 79868 173020 79932
rect 173084 79906 173116 79932
rect 173172 79906 173177 79962
rect 173084 79901 173177 79906
rect 173939 79962 174005 79967
rect 173939 79906 173944 79962
rect 174000 79930 174005 79962
rect 175963 79962 176029 79967
rect 175222 79930 175228 79932
rect 174000 79906 175228 79930
rect 173939 79901 175228 79906
rect 173084 79870 173128 79901
rect 173942 79870 175228 79901
rect 173084 79868 173090 79870
rect 175222 79868 175228 79870
rect 175292 79868 175298 79932
rect 175963 79906 175968 79962
rect 176024 79906 176029 79962
rect 175963 79901 176029 79906
rect 176331 79962 176397 79967
rect 176331 79906 176336 79962
rect 176392 79930 176397 79962
rect 177941 79930 178007 79933
rect 176392 79928 178007 79930
rect 176392 79906 177946 79928
rect 176331 79901 177946 79906
rect 172470 79792 172579 79797
rect 172470 79736 172518 79792
rect 172574 79736 172579 79792
rect 172470 79734 172579 79736
rect 172654 79794 172714 79867
rect 173065 79794 173131 79797
rect 174813 79796 174879 79797
rect 174813 79794 174860 79796
rect 172654 79792 173131 79794
rect 172654 79736 173070 79792
rect 173126 79736 173131 79792
rect 172654 79734 173131 79736
rect 174768 79792 174860 79794
rect 174768 79736 174818 79792
rect 174768 79734 174860 79736
rect 172513 79731 172579 79734
rect 173065 79731 173131 79734
rect 174813 79732 174860 79734
rect 174924 79732 174930 79796
rect 175966 79794 176026 79901
rect 176334 79872 177946 79901
rect 178002 79872 178007 79928
rect 176334 79870 178007 79872
rect 177941 79867 178007 79870
rect 180750 79870 186330 79930
rect 176745 79794 176811 79797
rect 177251 79796 177317 79797
rect 177246 79794 177252 79796
rect 175966 79792 176811 79794
rect 175966 79736 176750 79792
rect 176806 79736 176811 79792
rect 175966 79734 176811 79736
rect 177160 79734 177252 79794
rect 174813 79731 174879 79732
rect 176745 79731 176811 79734
rect 177246 79732 177252 79734
rect 177316 79732 177322 79796
rect 177251 79731 177317 79732
rect 180750 79658 180810 79870
rect 171918 79598 180810 79658
rect 166533 79595 166599 79596
rect 168741 79595 168807 79598
rect 171225 79595 171291 79598
rect 160369 79522 160435 79525
rect 155174 79520 160435 79522
rect 155174 79464 160374 79520
rect 160430 79464 160435 79520
rect 155174 79462 160435 79464
rect 154757 79459 154823 79462
rect 160369 79459 160435 79462
rect 162577 79522 162643 79525
rect 162710 79522 162716 79524
rect 162577 79520 162716 79522
rect 162577 79464 162582 79520
rect 162638 79464 162716 79520
rect 162577 79462 162716 79464
rect 162577 79459 162643 79462
rect 162710 79460 162716 79462
rect 162780 79460 162786 79524
rect 176694 79522 176700 79524
rect 165432 79462 176700 79522
rect 159633 79386 159699 79389
rect 165432 79386 165492 79462
rect 176694 79460 176700 79462
rect 176764 79460 176770 79524
rect 174721 79388 174787 79389
rect 174670 79386 174676 79388
rect 159633 79384 165492 79386
rect 159633 79328 159638 79384
rect 159694 79328 165492 79384
rect 159633 79326 165492 79328
rect 174630 79326 174676 79386
rect 174740 79384 174787 79388
rect 174782 79328 174787 79384
rect 159633 79323 159699 79326
rect 174670 79324 174676 79326
rect 174740 79324 174787 79328
rect 174721 79323 174787 79324
rect 175365 79386 175431 79389
rect 176510 79386 176516 79388
rect 175365 79384 176516 79386
rect 175365 79328 175370 79384
rect 175426 79328 176516 79384
rect 175365 79326 176516 79328
rect 175365 79323 175431 79326
rect 176510 79324 176516 79326
rect 176580 79324 176586 79388
rect 186270 79386 186330 79870
rect 212809 79386 212875 79389
rect 186270 79384 212875 79386
rect 186270 79328 212814 79384
rect 212870 79328 212875 79384
rect 186270 79326 212875 79328
rect 212809 79323 212875 79326
rect 168373 79250 168439 79253
rect 151632 79248 168439 79250
rect 151632 79192 168378 79248
rect 168434 79192 168439 79248
rect 151632 79190 168439 79192
rect 139301 79187 139367 79188
rect 140773 79187 140839 79190
rect 141233 79187 141299 79190
rect 168373 79187 168439 79190
rect 171225 79250 171291 79253
rect 184790 79250 184796 79252
rect 171225 79248 184796 79250
rect 171225 79192 171230 79248
rect 171286 79192 184796 79248
rect 171225 79190 184796 79192
rect 171225 79187 171291 79190
rect 184790 79188 184796 79190
rect 184860 79188 184866 79252
rect 139894 79052 139900 79116
rect 139964 79114 139970 79116
rect 142337 79114 142403 79117
rect 139964 79112 142403 79114
rect 139964 79056 142342 79112
rect 142398 79056 142403 79112
rect 139964 79054 142403 79056
rect 139964 79052 139970 79054
rect 142337 79051 142403 79054
rect 142654 79052 142660 79116
rect 142724 79114 142730 79116
rect 142797 79114 142863 79117
rect 142724 79112 142863 79114
rect 142724 79056 142802 79112
rect 142858 79056 142863 79112
rect 142724 79054 142863 79056
rect 142724 79052 142730 79054
rect 142797 79051 142863 79054
rect 156873 79114 156939 79117
rect 186313 79114 186379 79117
rect 156873 79112 186379 79114
rect 156873 79056 156878 79112
rect 156934 79056 186318 79112
rect 186374 79056 186379 79112
rect 156873 79054 186379 79056
rect 156873 79051 156939 79054
rect 186313 79051 186379 79054
rect 153745 78978 153811 78981
rect 167821 78980 167887 78981
rect 168281 78980 168347 78981
rect 170857 78980 170923 78981
rect 167821 78978 167868 78980
rect 137970 78976 153811 78978
rect 137970 78920 153750 78976
rect 153806 78920 153811 78976
rect 137970 78918 153811 78920
rect 167776 78976 167868 78978
rect 167776 78920 167826 78976
rect 167776 78918 167868 78920
rect 102869 78915 102935 78918
rect 137461 78915 137527 78918
rect 153745 78915 153811 78918
rect 167821 78916 167868 78918
rect 167932 78916 167938 78980
rect 168230 78916 168236 78980
rect 168300 78978 168347 78980
rect 168300 78976 168392 78978
rect 168342 78920 168392 78976
rect 168300 78918 168392 78920
rect 168300 78916 168347 78918
rect 170806 78916 170812 78980
rect 170876 78978 170923 78980
rect 172697 78978 172763 78981
rect 214373 78978 214439 78981
rect 170876 78976 170968 78978
rect 170918 78920 170968 78976
rect 170876 78918 170968 78920
rect 172697 78976 214439 78978
rect 172697 78920 172702 78976
rect 172758 78920 214378 78976
rect 214434 78920 214439 78976
rect 172697 78918 214439 78920
rect 170876 78916 170923 78918
rect 167821 78915 167887 78916
rect 168281 78915 168347 78916
rect 170857 78915 170923 78916
rect 172697 78915 172763 78918
rect 214373 78915 214439 78918
rect 109493 78842 109559 78845
rect 144361 78842 144427 78845
rect 109493 78840 144427 78842
rect 109493 78784 109498 78840
rect 109554 78784 144366 78840
rect 144422 78784 144427 78840
rect 109493 78782 144427 78784
rect 109493 78779 109559 78782
rect 144361 78779 144427 78782
rect 167126 78780 167132 78844
rect 167196 78842 167202 78844
rect 167862 78842 167868 78844
rect 167196 78782 167868 78842
rect 167196 78780 167202 78782
rect 167862 78780 167868 78782
rect 167932 78780 167938 78844
rect 169477 78842 169543 78845
rect 214465 78842 214531 78845
rect 169477 78840 214531 78842
rect 169477 78784 169482 78840
rect 169538 78784 214470 78840
rect 214526 78784 214531 78840
rect 169477 78782 214531 78784
rect 169477 78779 169543 78782
rect 214465 78779 214531 78782
rect 99230 78644 99236 78708
rect 99300 78706 99306 78708
rect 154062 78706 154068 78708
rect 99300 78646 154068 78706
rect 99300 78644 99306 78646
rect 154062 78644 154068 78646
rect 154132 78644 154138 78708
rect 156086 78644 156092 78708
rect 156156 78706 156162 78708
rect 156413 78706 156479 78709
rect 156156 78704 156479 78706
rect 156156 78648 156418 78704
rect 156474 78648 156479 78704
rect 156156 78646 156479 78648
rect 156156 78644 156162 78646
rect 156413 78643 156479 78646
rect 161105 78706 161171 78709
rect 161238 78706 161244 78708
rect 161105 78704 161244 78706
rect 161105 78648 161110 78704
rect 161166 78648 161244 78704
rect 161105 78646 161244 78648
rect 161105 78643 161171 78646
rect 161238 78644 161244 78646
rect 161308 78644 161314 78708
rect 163446 78644 163452 78708
rect 163516 78706 163522 78708
rect 217317 78706 217383 78709
rect 163516 78704 217383 78706
rect 163516 78648 217322 78704
rect 217378 78648 217383 78704
rect 163516 78646 217383 78648
rect 163516 78644 163522 78646
rect 217317 78643 217383 78646
rect 119286 78508 119292 78572
rect 119356 78570 119362 78572
rect 119981 78570 120047 78573
rect 122281 78572 122347 78573
rect 122230 78570 122236 78572
rect 119356 78568 120047 78570
rect 119356 78512 119986 78568
rect 120042 78512 120047 78568
rect 119356 78510 120047 78512
rect 122190 78510 122236 78570
rect 122300 78568 122347 78572
rect 128445 78570 128511 78573
rect 122342 78512 122347 78568
rect 119356 78508 119362 78510
rect 119981 78507 120047 78510
rect 122230 78508 122236 78510
rect 122300 78508 122347 78512
rect 122281 78507 122347 78508
rect 122790 78568 128511 78570
rect 122790 78512 128450 78568
rect 128506 78512 128511 78568
rect 122790 78510 128511 78512
rect 100334 78372 100340 78436
rect 100404 78434 100410 78436
rect 122790 78434 122850 78510
rect 128445 78507 128511 78510
rect 134609 78570 134675 78573
rect 134926 78570 134932 78572
rect 134609 78568 134932 78570
rect 134609 78512 134614 78568
rect 134670 78512 134932 78568
rect 134609 78510 134932 78512
rect 134609 78507 134675 78510
rect 134926 78508 134932 78510
rect 134996 78508 135002 78572
rect 140446 78508 140452 78572
rect 140516 78570 140522 78572
rect 143441 78570 143507 78573
rect 140516 78568 143507 78570
rect 140516 78512 143446 78568
rect 143502 78512 143507 78568
rect 140516 78510 143507 78512
rect 140516 78508 140522 78510
rect 143441 78507 143507 78510
rect 156597 78572 156663 78573
rect 156597 78568 156644 78572
rect 156708 78570 156714 78572
rect 156597 78512 156602 78568
rect 156597 78508 156644 78512
rect 156708 78510 156754 78570
rect 156708 78508 156714 78510
rect 159582 78508 159588 78572
rect 159652 78570 159658 78572
rect 162669 78570 162735 78573
rect 159652 78568 162735 78570
rect 159652 78512 162674 78568
rect 162730 78512 162735 78568
rect 159652 78510 162735 78512
rect 159652 78508 159658 78510
rect 156597 78507 156663 78508
rect 162669 78507 162735 78510
rect 164601 78570 164667 78573
rect 164918 78570 164924 78572
rect 164601 78568 164924 78570
rect 164601 78512 164606 78568
rect 164662 78512 164924 78568
rect 164601 78510 164924 78512
rect 164601 78507 164667 78510
rect 164918 78508 164924 78510
rect 164988 78508 164994 78572
rect 165981 78570 166047 78573
rect 171726 78570 171732 78572
rect 165981 78568 171732 78570
rect 165981 78512 165986 78568
rect 166042 78512 171732 78568
rect 165981 78510 171732 78512
rect 165981 78507 166047 78510
rect 171726 78508 171732 78510
rect 171796 78508 171802 78572
rect 177573 78570 177639 78573
rect 213085 78570 213151 78573
rect 177573 78568 213151 78570
rect 177573 78512 177578 78568
rect 177634 78512 213090 78568
rect 213146 78512 213151 78568
rect 177573 78510 213151 78512
rect 177573 78507 177639 78510
rect 213085 78507 213151 78510
rect 100404 78374 122850 78434
rect 100404 78372 100410 78374
rect 123886 78372 123892 78436
rect 123956 78434 123962 78436
rect 124581 78434 124647 78437
rect 123956 78432 124647 78434
rect 123956 78376 124586 78432
rect 124642 78376 124647 78432
rect 123956 78374 124647 78376
rect 123956 78372 123962 78374
rect 124581 78371 124647 78374
rect 135069 78434 135135 78437
rect 135662 78434 135668 78436
rect 135069 78432 135668 78434
rect 135069 78376 135074 78432
rect 135130 78376 135668 78432
rect 135069 78374 135668 78376
rect 135069 78371 135135 78374
rect 135662 78372 135668 78374
rect 135732 78372 135738 78436
rect 142102 78372 142108 78436
rect 142172 78434 142178 78436
rect 143073 78434 143139 78437
rect 142172 78432 143139 78434
rect 142172 78376 143078 78432
rect 143134 78376 143139 78432
rect 142172 78374 143139 78376
rect 142172 78372 142178 78374
rect 143073 78371 143139 78374
rect 145005 78434 145071 78437
rect 149278 78434 149284 78436
rect 145005 78432 149284 78434
rect 145005 78376 145010 78432
rect 145066 78376 149284 78432
rect 145005 78374 149284 78376
rect 145005 78371 145071 78374
rect 149278 78372 149284 78374
rect 149348 78372 149354 78436
rect 163865 78434 163931 78437
rect 175089 78434 175155 78437
rect 183921 78434 183987 78437
rect 184197 78434 184263 78437
rect 163865 78432 168298 78434
rect 163865 78376 163870 78432
rect 163926 78376 168298 78432
rect 163865 78374 168298 78376
rect 163865 78371 163931 78374
rect 100518 78236 100524 78300
rect 100588 78298 100594 78300
rect 128629 78298 128695 78301
rect 100588 78296 128695 78298
rect 100588 78240 128634 78296
rect 128690 78240 128695 78296
rect 100588 78238 128695 78240
rect 100588 78236 100594 78238
rect 128629 78235 128695 78238
rect 147990 78236 147996 78300
rect 148060 78298 148066 78300
rect 148593 78298 148659 78301
rect 148060 78296 148659 78298
rect 148060 78240 148598 78296
rect 148654 78240 148659 78296
rect 148060 78238 148659 78240
rect 148060 78236 148066 78238
rect 148593 78235 148659 78238
rect 150934 78236 150940 78300
rect 151004 78298 151010 78300
rect 151169 78298 151235 78301
rect 151004 78296 151235 78298
rect 151004 78240 151174 78296
rect 151230 78240 151235 78296
rect 151004 78238 151235 78240
rect 151004 78236 151010 78238
rect 151169 78235 151235 78238
rect 157977 78298 158043 78301
rect 165838 78298 165844 78300
rect 157977 78296 165844 78298
rect 157977 78240 157982 78296
rect 158038 78240 165844 78296
rect 157977 78238 165844 78240
rect 157977 78235 158043 78238
rect 165838 78236 165844 78238
rect 165908 78236 165914 78300
rect 168238 78298 168298 78374
rect 175089 78432 184263 78434
rect 175089 78376 175094 78432
rect 175150 78376 183926 78432
rect 183982 78376 184202 78432
rect 184258 78376 184263 78432
rect 175089 78374 184263 78376
rect 175089 78371 175155 78374
rect 183921 78371 183987 78374
rect 184197 78371 184263 78374
rect 186313 78434 186379 78437
rect 186998 78434 187004 78436
rect 186313 78432 187004 78434
rect 186313 78376 186318 78432
rect 186374 78376 187004 78432
rect 186313 78374 187004 78376
rect 186313 78371 186379 78374
rect 186998 78372 187004 78374
rect 187068 78372 187074 78436
rect 195421 78298 195487 78301
rect 168238 78296 195487 78298
rect 168238 78240 195426 78296
rect 195482 78240 195487 78296
rect 168238 78238 195487 78240
rect 195421 78235 195487 78238
rect 124070 78100 124076 78164
rect 124140 78162 124146 78164
rect 134609 78162 134675 78165
rect 141233 78164 141299 78165
rect 124140 78160 134675 78162
rect 124140 78104 134614 78160
rect 134670 78104 134675 78160
rect 124140 78102 134675 78104
rect 124140 78100 124146 78102
rect 134609 78099 134675 78102
rect 141182 78100 141188 78164
rect 141252 78162 141299 78164
rect 144361 78162 144427 78165
rect 144494 78162 144500 78164
rect 141252 78160 141344 78162
rect 141294 78104 141344 78160
rect 141252 78102 141344 78104
rect 144361 78160 144500 78162
rect 144361 78104 144366 78160
rect 144422 78104 144500 78160
rect 144361 78102 144500 78104
rect 141252 78100 141299 78102
rect 141233 78099 141299 78100
rect 144361 78099 144427 78102
rect 144494 78100 144500 78102
rect 144564 78100 144570 78164
rect 150617 78162 150683 78165
rect 173065 78164 173131 78165
rect 161974 78162 161980 78164
rect 150617 78160 161980 78162
rect 150617 78104 150622 78160
rect 150678 78104 161980 78160
rect 150617 78102 161980 78104
rect 150617 78099 150683 78102
rect 161974 78100 161980 78102
rect 162044 78100 162050 78164
rect 173014 78100 173020 78164
rect 173084 78162 173131 78164
rect 174721 78162 174787 78165
rect 182173 78162 182239 78165
rect 189206 78162 189212 78164
rect 173084 78160 173176 78162
rect 173126 78104 173176 78160
rect 173084 78102 173176 78104
rect 174721 78160 180810 78162
rect 174721 78104 174726 78160
rect 174782 78104 180810 78160
rect 174721 78102 180810 78104
rect 173084 78100 173131 78102
rect 173065 78099 173131 78100
rect 174721 78099 174787 78102
rect 121126 77964 121132 78028
rect 121196 78026 121202 78028
rect 134885 78026 134951 78029
rect 121196 78024 134951 78026
rect 121196 77968 134890 78024
rect 134946 77968 134951 78024
rect 121196 77966 134951 77968
rect 121196 77964 121202 77966
rect 134885 77963 134951 77966
rect 139342 77964 139348 78028
rect 139412 78026 139418 78028
rect 146017 78026 146083 78029
rect 139412 78024 146083 78026
rect 139412 77968 146022 78024
rect 146078 77968 146083 78024
rect 139412 77966 146083 77968
rect 139412 77964 139418 77966
rect 146017 77963 146083 77966
rect 146702 77964 146708 78028
rect 146772 78026 146778 78028
rect 147305 78026 147371 78029
rect 146772 78024 147371 78026
rect 146772 77968 147310 78024
rect 147366 77968 147371 78024
rect 146772 77966 147371 77968
rect 146772 77964 146778 77966
rect 147305 77963 147371 77966
rect 149278 77964 149284 78028
rect 149348 78026 149354 78028
rect 149421 78026 149487 78029
rect 149348 78024 149487 78026
rect 149348 77968 149426 78024
rect 149482 77968 149487 78024
rect 149348 77966 149487 77968
rect 149348 77964 149354 77966
rect 149421 77963 149487 77966
rect 149646 77964 149652 78028
rect 149716 78026 149722 78028
rect 150249 78026 150315 78029
rect 149716 78024 150315 78026
rect 149716 77968 150254 78024
rect 150310 77968 150315 78024
rect 149716 77966 150315 77968
rect 149716 77964 149722 77966
rect 150249 77963 150315 77966
rect 153285 78026 153351 78029
rect 153694 78026 153700 78028
rect 153285 78024 153700 78026
rect 153285 77968 153290 78024
rect 153346 77968 153700 78024
rect 153285 77966 153700 77968
rect 153285 77963 153351 77966
rect 153694 77964 153700 77966
rect 153764 77964 153770 78028
rect 165797 78026 165863 78029
rect 175038 78026 175044 78028
rect 165797 78024 175044 78026
rect 165797 77968 165802 78024
rect 165858 77968 175044 78024
rect 165797 77966 175044 77968
rect 165797 77963 165863 77966
rect 175038 77964 175044 77966
rect 175108 77964 175114 78028
rect 180750 78026 180810 78102
rect 182173 78160 189212 78162
rect 182173 78104 182178 78160
rect 182234 78104 189212 78160
rect 182173 78102 189212 78104
rect 182173 78099 182239 78102
rect 189206 78100 189212 78102
rect 189276 78100 189282 78164
rect 189022 78026 189028 78028
rect 180750 77966 189028 78026
rect 189022 77964 189028 77966
rect 189092 77964 189098 78028
rect 140037 77890 140103 77893
rect 131070 77888 140103 77890
rect 131070 77832 140042 77888
rect 140098 77832 140103 77888
rect 131070 77830 140103 77832
rect 107142 77692 107148 77756
rect 107212 77754 107218 77756
rect 131070 77754 131130 77830
rect 140037 77827 140103 77830
rect 143574 77828 143580 77892
rect 143644 77890 143650 77892
rect 144453 77890 144519 77893
rect 143644 77888 144519 77890
rect 143644 77832 144458 77888
rect 144514 77832 144519 77888
rect 143644 77830 144519 77832
rect 143644 77828 143650 77830
rect 144453 77827 144519 77830
rect 152774 77828 152780 77892
rect 152844 77890 152850 77892
rect 170806 77890 170812 77892
rect 152844 77830 170812 77890
rect 152844 77828 152850 77830
rect 170806 77828 170812 77830
rect 170876 77828 170882 77892
rect 179965 77890 180031 77893
rect 215937 77890 216003 77893
rect 179965 77888 216003 77890
rect 179965 77832 179970 77888
rect 180026 77832 215942 77888
rect 215998 77832 216003 77888
rect 179965 77830 216003 77832
rect 179965 77827 180031 77830
rect 215937 77827 216003 77830
rect 107212 77694 131130 77754
rect 107212 77692 107218 77694
rect 135846 77692 135852 77756
rect 135916 77754 135922 77756
rect 137093 77754 137159 77757
rect 135916 77752 137159 77754
rect 135916 77696 137098 77752
rect 137154 77696 137159 77752
rect 135916 77694 137159 77696
rect 135916 77692 135922 77694
rect 137093 77691 137159 77694
rect 144126 77692 144132 77756
rect 144196 77754 144202 77756
rect 151721 77754 151787 77757
rect 144196 77752 151787 77754
rect 144196 77696 151726 77752
rect 151782 77696 151787 77752
rect 144196 77694 151787 77696
rect 144196 77692 144202 77694
rect 151721 77691 151787 77694
rect 179045 77754 179111 77757
rect 211429 77754 211495 77757
rect 179045 77752 211495 77754
rect 179045 77696 179050 77752
rect 179106 77696 211434 77752
rect 211490 77696 211495 77752
rect 179045 77694 211495 77696
rect 179045 77691 179111 77694
rect 211429 77691 211495 77694
rect 120942 77556 120948 77620
rect 121012 77618 121018 77620
rect 137737 77618 137803 77621
rect 121012 77616 137803 77618
rect 121012 77560 137742 77616
rect 137798 77560 137803 77616
rect 121012 77558 137803 77560
rect 121012 77556 121018 77558
rect 137737 77555 137803 77558
rect 138238 77556 138244 77620
rect 138308 77618 138314 77620
rect 138749 77618 138815 77621
rect 138308 77616 138815 77618
rect 138308 77560 138754 77616
rect 138810 77560 138815 77616
rect 138308 77558 138815 77560
rect 138308 77556 138314 77558
rect 138749 77555 138815 77558
rect 151537 77618 151603 77621
rect 162894 77618 162900 77620
rect 151537 77616 162900 77618
rect 151537 77560 151542 77616
rect 151598 77560 162900 77616
rect 151537 77558 162900 77560
rect 151537 77555 151603 77558
rect 162894 77556 162900 77558
rect 162964 77556 162970 77620
rect 101673 77210 101739 77213
rect 135713 77210 135779 77213
rect 101673 77208 135779 77210
rect 101673 77152 101678 77208
rect 101734 77152 135718 77208
rect 135774 77152 135779 77208
rect 101673 77150 135779 77152
rect 101673 77147 101739 77150
rect 135713 77147 135779 77150
rect 154665 77210 154731 77213
rect 160686 77210 160692 77212
rect 154665 77208 160692 77210
rect 154665 77152 154670 77208
rect 154726 77152 160692 77208
rect 154665 77150 160692 77152
rect 154665 77147 154731 77150
rect 160686 77148 160692 77150
rect 160756 77148 160762 77212
rect 162025 77210 162091 77213
rect 189625 77210 189691 77213
rect 162025 77208 189691 77210
rect 162025 77152 162030 77208
rect 162086 77152 189630 77208
rect 189686 77152 189691 77208
rect 162025 77150 189691 77152
rect 162025 77147 162091 77150
rect 189625 77147 189691 77150
rect 159817 77074 159883 77077
rect 217225 77074 217291 77077
rect 159817 77072 217291 77074
rect 159817 77016 159822 77072
rect 159878 77016 217230 77072
rect 217286 77016 217291 77072
rect 159817 77014 217291 77016
rect 159817 77011 159883 77014
rect 217225 77011 217291 77014
rect 108205 76938 108271 76941
rect 138657 76938 138723 76941
rect 108205 76936 138723 76938
rect 108205 76880 108210 76936
rect 108266 76880 138662 76936
rect 138718 76880 138723 76936
rect 108205 76878 138723 76880
rect 108205 76875 108271 76878
rect 138657 76875 138723 76878
rect 170806 76876 170812 76940
rect 170876 76938 170882 76940
rect 218513 76938 218579 76941
rect 170876 76936 218579 76938
rect 170876 76880 218518 76936
rect 218574 76880 218579 76936
rect 170876 76878 218579 76880
rect 170876 76876 170882 76878
rect 218513 76875 218579 76878
rect 580625 76938 580691 76941
rect 583520 76938 584960 77028
rect 580625 76936 584960 76938
rect 580625 76880 580630 76936
rect 580686 76880 584960 76936
rect 580625 76878 584960 76880
rect 580625 76875 580691 76878
rect 108430 76740 108436 76804
rect 108500 76802 108506 76804
rect 136633 76802 136699 76805
rect 140221 76804 140287 76805
rect 140221 76802 140268 76804
rect 108500 76800 136699 76802
rect 108500 76744 136638 76800
rect 136694 76744 136699 76800
rect 108500 76742 136699 76744
rect 140176 76800 140268 76802
rect 140176 76744 140226 76800
rect 140176 76742 140268 76744
rect 108500 76740 108506 76742
rect 136633 76739 136699 76742
rect 140221 76740 140268 76742
rect 140332 76740 140338 76804
rect 177297 76802 177363 76805
rect 209957 76802 210023 76805
rect 210366 76802 210372 76804
rect 177297 76800 200130 76802
rect 177297 76744 177302 76800
rect 177358 76744 200130 76800
rect 177297 76742 200130 76744
rect 140221 76739 140287 76740
rect 177297 76739 177363 76742
rect 119838 76604 119844 76668
rect 119908 76666 119914 76668
rect 147949 76666 148015 76669
rect 119908 76664 148015 76666
rect 119908 76608 147954 76664
rect 148010 76608 148015 76664
rect 119908 76606 148015 76608
rect 119908 76604 119914 76606
rect 147949 76603 148015 76606
rect 158069 76668 158135 76669
rect 158069 76664 158116 76668
rect 158180 76666 158186 76668
rect 158069 76608 158074 76664
rect 158069 76604 158116 76608
rect 158180 76606 158226 76666
rect 158180 76604 158186 76606
rect 158294 76604 158300 76668
rect 158364 76666 158370 76668
rect 158437 76666 158503 76669
rect 158364 76664 158503 76666
rect 158364 76608 158442 76664
rect 158498 76608 158503 76664
rect 158364 76606 158503 76608
rect 158364 76604 158370 76606
rect 158069 76603 158135 76604
rect 158437 76603 158503 76606
rect 164969 76666 165035 76669
rect 198774 76666 198780 76668
rect 164969 76664 198780 76666
rect 164969 76608 164974 76664
rect 165030 76608 198780 76664
rect 164969 76606 198780 76608
rect 164969 76603 165035 76606
rect 198774 76604 198780 76606
rect 198844 76604 198850 76668
rect 200070 76666 200130 76742
rect 209957 76800 210372 76802
rect 209957 76744 209962 76800
rect 210018 76744 210372 76800
rect 209957 76742 210372 76744
rect 209957 76739 210023 76742
rect 210366 76740 210372 76742
rect 210436 76740 210442 76804
rect 583520 76788 584960 76878
rect 211102 76666 211108 76668
rect 200070 76606 211108 76666
rect 211102 76604 211108 76606
rect 211172 76604 211178 76668
rect 115422 76468 115428 76532
rect 115492 76530 115498 76532
rect 144545 76530 144611 76533
rect 115492 76528 144611 76530
rect 115492 76472 144550 76528
rect 144606 76472 144611 76528
rect 115492 76470 144611 76472
rect 115492 76468 115498 76470
rect 144545 76467 144611 76470
rect 164877 76530 164943 76533
rect 174629 76530 174695 76533
rect 164877 76528 174695 76530
rect 164877 76472 164882 76528
rect 164938 76472 174634 76528
rect 174690 76472 174695 76528
rect 164877 76470 174695 76472
rect 164877 76467 164943 76470
rect 174629 76467 174695 76470
rect 177941 76530 178007 76533
rect 200389 76530 200455 76533
rect 177941 76528 200455 76530
rect 177941 76472 177946 76528
rect 178002 76472 200394 76528
rect 200450 76472 200455 76528
rect 177941 76470 200455 76472
rect 177941 76467 178007 76470
rect 200389 76467 200455 76470
rect 139577 76394 139643 76397
rect 140078 76394 140084 76396
rect 139577 76392 140084 76394
rect -960 76258 480 76348
rect 139577 76336 139582 76392
rect 139638 76336 140084 76392
rect 139577 76334 140084 76336
rect 139577 76331 139643 76334
rect 140078 76332 140084 76334
rect 140148 76332 140154 76396
rect 155401 76394 155467 76397
rect 215385 76394 215451 76397
rect 155401 76392 215451 76394
rect 155401 76336 155406 76392
rect 155462 76336 215390 76392
rect 215446 76336 215451 76392
rect 155401 76334 215451 76336
rect 155401 76331 155467 76334
rect 215385 76331 215451 76334
rect 2773 76258 2839 76261
rect -960 76256 2839 76258
rect -960 76200 2778 76256
rect 2834 76200 2839 76256
rect -960 76198 2839 76200
rect -960 76108 480 76198
rect 2773 76195 2839 76198
rect 116393 76258 116459 76261
rect 148542 76258 148548 76260
rect 116393 76256 148548 76258
rect 116393 76200 116398 76256
rect 116454 76200 148548 76256
rect 116393 76198 148548 76200
rect 116393 76195 116459 76198
rect 148542 76196 148548 76198
rect 148612 76196 148618 76260
rect 136081 76122 136147 76125
rect 136214 76122 136220 76124
rect 136081 76120 136220 76122
rect 136081 76064 136086 76120
rect 136142 76064 136220 76120
rect 136081 76062 136220 76064
rect 136081 76059 136147 76062
rect 136214 76060 136220 76062
rect 136284 76060 136290 76124
rect 169753 76122 169819 76125
rect 170622 76122 170628 76124
rect 169753 76120 170628 76122
rect 169753 76064 169758 76120
rect 169814 76064 170628 76120
rect 169753 76062 170628 76064
rect 169753 76059 169819 76062
rect 170622 76060 170628 76062
rect 170692 76060 170698 76124
rect 132585 75986 132651 75989
rect 136357 75988 136423 75989
rect 158805 75988 158871 75989
rect 160461 75988 160527 75989
rect 170029 75988 170095 75989
rect 133086 75986 133092 75988
rect 132585 75984 133092 75986
rect 132585 75928 132590 75984
rect 132646 75928 133092 75984
rect 132585 75926 133092 75928
rect 132585 75923 132651 75926
rect 133086 75924 133092 75926
rect 133156 75924 133162 75988
rect 136357 75986 136404 75988
rect 136312 75984 136404 75986
rect 136312 75928 136362 75984
rect 136312 75926 136404 75928
rect 136357 75924 136404 75926
rect 136468 75924 136474 75988
rect 158805 75986 158852 75988
rect 158760 75984 158852 75986
rect 158760 75928 158810 75984
rect 158760 75926 158852 75928
rect 158805 75924 158852 75926
rect 158916 75924 158922 75988
rect 160461 75986 160508 75988
rect 160416 75984 160508 75986
rect 160416 75928 160466 75984
rect 160416 75926 160508 75928
rect 160461 75924 160508 75926
rect 160572 75924 160578 75988
rect 170029 75986 170076 75988
rect 169984 75984 170076 75986
rect 169984 75928 170034 75984
rect 169984 75926 170076 75928
rect 170029 75924 170076 75926
rect 170140 75924 170146 75988
rect 171961 75986 172027 75989
rect 172278 75986 172284 75988
rect 171961 75984 172284 75986
rect 171961 75928 171966 75984
rect 172022 75928 172284 75984
rect 171961 75926 172284 75928
rect 136357 75923 136423 75924
rect 158805 75923 158871 75924
rect 160461 75923 160527 75924
rect 170029 75923 170095 75924
rect 171961 75923 172027 75926
rect 172278 75924 172284 75926
rect 172348 75924 172354 75988
rect 119797 75850 119863 75853
rect 145649 75850 145715 75853
rect 119797 75848 145715 75850
rect 119797 75792 119802 75848
rect 119858 75792 145654 75848
rect 145710 75792 145715 75848
rect 119797 75790 145715 75792
rect 119797 75787 119863 75790
rect 145649 75787 145715 75790
rect 160093 75850 160159 75853
rect 163446 75850 163452 75852
rect 160093 75848 163452 75850
rect 160093 75792 160098 75848
rect 160154 75792 163452 75848
rect 160093 75790 163452 75792
rect 160093 75787 160159 75790
rect 163446 75788 163452 75790
rect 163516 75788 163522 75852
rect 176009 75850 176075 75853
rect 209037 75850 209103 75853
rect 176009 75848 209103 75850
rect 176009 75792 176014 75848
rect 176070 75792 209042 75848
rect 209098 75792 209103 75848
rect 176009 75790 209103 75792
rect 176009 75787 176075 75790
rect 209037 75787 209103 75790
rect 97073 75714 97139 75717
rect 143942 75714 143948 75716
rect 97073 75712 143948 75714
rect 97073 75656 97078 75712
rect 97134 75656 143948 75712
rect 97073 75654 143948 75656
rect 97073 75651 97139 75654
rect 143942 75652 143948 75654
rect 144012 75652 144018 75716
rect 173801 75714 173867 75717
rect 214005 75714 214071 75717
rect 173801 75712 214071 75714
rect 173801 75656 173806 75712
rect 173862 75656 214010 75712
rect 214066 75656 214071 75712
rect 173801 75654 214071 75656
rect 173801 75651 173867 75654
rect 214005 75651 214071 75654
rect 114921 75578 114987 75581
rect 148409 75578 148475 75581
rect 114921 75576 148475 75578
rect 114921 75520 114926 75576
rect 114982 75520 148414 75576
rect 148470 75520 148475 75576
rect 114921 75518 148475 75520
rect 114921 75515 114987 75518
rect 148409 75515 148475 75518
rect 173157 75578 173223 75581
rect 212625 75578 212691 75581
rect 173157 75576 212691 75578
rect 173157 75520 173162 75576
rect 173218 75520 212630 75576
rect 212686 75520 212691 75576
rect 173157 75518 212691 75520
rect 173157 75515 173223 75518
rect 212625 75515 212691 75518
rect 109401 75442 109467 75445
rect 140630 75442 140636 75444
rect 109401 75440 140636 75442
rect 109401 75384 109406 75440
rect 109462 75384 140636 75440
rect 109401 75382 140636 75384
rect 109401 75379 109467 75382
rect 140630 75380 140636 75382
rect 140700 75380 140706 75444
rect 178953 75442 179019 75445
rect 214046 75442 214052 75444
rect 178953 75440 214052 75442
rect 178953 75384 178958 75440
rect 179014 75384 214052 75440
rect 178953 75382 214052 75384
rect 178953 75379 179019 75382
rect 214046 75380 214052 75382
rect 214116 75380 214122 75444
rect 117078 75244 117084 75308
rect 117148 75306 117154 75308
rect 146702 75306 146708 75308
rect 117148 75246 146708 75306
rect 117148 75244 117154 75246
rect 146702 75244 146708 75246
rect 146772 75244 146778 75308
rect 176193 75306 176259 75309
rect 210325 75306 210391 75309
rect 176193 75304 210391 75306
rect 176193 75248 176198 75304
rect 176254 75248 210330 75304
rect 210386 75248 210391 75304
rect 176193 75246 210391 75248
rect 176193 75243 176259 75246
rect 210325 75243 210391 75246
rect 114134 75108 114140 75172
rect 114204 75170 114210 75172
rect 136725 75170 136791 75173
rect 114204 75168 136791 75170
rect 114204 75112 136730 75168
rect 136786 75112 136791 75168
rect 114204 75110 136791 75112
rect 114204 75108 114210 75110
rect 136725 75107 136791 75110
rect 96981 75034 97047 75037
rect 145189 75034 145255 75037
rect 96981 75032 145255 75034
rect 96981 74976 96986 75032
rect 97042 74976 145194 75032
rect 145250 74976 145255 75032
rect 96981 74974 145255 74976
rect 96981 74971 97047 74974
rect 145189 74971 145255 74974
rect 153561 75034 153627 75037
rect 199193 75034 199259 75037
rect 153561 75032 199259 75034
rect 153561 74976 153566 75032
rect 153622 74976 199198 75032
rect 199254 74976 199259 75032
rect 153561 74974 199259 74976
rect 153561 74971 153627 74974
rect 199193 74971 199259 74974
rect 128445 74490 128511 74493
rect 139393 74490 139459 74493
rect 128445 74488 139459 74490
rect 128445 74432 128450 74488
rect 128506 74432 139398 74488
rect 139454 74432 139459 74488
rect 128445 74430 139459 74432
rect 128445 74427 128511 74430
rect 139393 74427 139459 74430
rect 162342 74428 162348 74492
rect 162412 74490 162418 74492
rect 188429 74490 188495 74493
rect 162412 74488 188495 74490
rect 162412 74432 188434 74488
rect 188490 74432 188495 74488
rect 162412 74430 188495 74432
rect 162412 74428 162418 74430
rect 188429 74427 188495 74430
rect 118366 74292 118372 74356
rect 118436 74354 118442 74356
rect 152590 74354 152596 74356
rect 118436 74294 152596 74354
rect 118436 74292 118442 74294
rect 152590 74292 152596 74294
rect 152660 74292 152666 74356
rect 174670 74292 174676 74356
rect 174740 74354 174746 74356
rect 181437 74354 181503 74357
rect 174740 74352 181503 74354
rect 174740 74296 181442 74352
rect 181498 74296 181503 74352
rect 174740 74294 181503 74296
rect 174740 74292 174746 74294
rect 181437 74291 181503 74294
rect 99189 74218 99255 74221
rect 133505 74218 133571 74221
rect 99189 74216 133571 74218
rect 99189 74160 99194 74216
rect 99250 74160 133510 74216
rect 133566 74160 133571 74216
rect 99189 74158 133571 74160
rect 99189 74155 99255 74158
rect 133505 74155 133571 74158
rect 156086 74156 156092 74220
rect 156156 74218 156162 74220
rect 190494 74218 190500 74220
rect 156156 74158 190500 74218
rect 156156 74156 156162 74158
rect 190494 74156 190500 74158
rect 190564 74156 190570 74220
rect 118182 74020 118188 74084
rect 118252 74082 118258 74084
rect 150893 74082 150959 74085
rect 118252 74080 150959 74082
rect 118252 74024 150898 74080
rect 150954 74024 150959 74080
rect 118252 74022 150959 74024
rect 118252 74020 118258 74022
rect 150893 74019 150959 74022
rect 163630 74020 163636 74084
rect 163700 74082 163706 74084
rect 196198 74082 196204 74084
rect 163700 74022 196204 74082
rect 163700 74020 163706 74022
rect 196198 74020 196204 74022
rect 196268 74020 196274 74084
rect 108665 73946 108731 73949
rect 140446 73946 140452 73948
rect 108665 73944 140452 73946
rect 108665 73888 108670 73944
rect 108726 73888 140452 73944
rect 108665 73886 140452 73888
rect 108665 73883 108731 73886
rect 140446 73884 140452 73886
rect 140516 73884 140522 73948
rect 171726 73884 171732 73948
rect 171796 73946 171802 73948
rect 200573 73946 200639 73949
rect 171796 73944 200639 73946
rect 171796 73888 200578 73944
rect 200634 73888 200639 73944
rect 171796 73886 200639 73888
rect 171796 73884 171802 73886
rect 200573 73883 200639 73886
rect 115606 73748 115612 73812
rect 115676 73810 115682 73812
rect 146937 73810 147003 73813
rect 115676 73808 147003 73810
rect 115676 73752 146942 73808
rect 146998 73752 147003 73808
rect 115676 73750 147003 73752
rect 115676 73748 115682 73750
rect 146937 73747 147003 73750
rect 160001 73810 160067 73813
rect 193622 73810 193628 73812
rect 160001 73808 193628 73810
rect 160001 73752 160006 73808
rect 160062 73752 193628 73808
rect 160001 73750 193628 73752
rect 160001 73747 160067 73750
rect 193622 73748 193628 73750
rect 193692 73748 193698 73812
rect 113030 73612 113036 73676
rect 113100 73674 113106 73676
rect 153101 73674 153167 73677
rect 113100 73672 153167 73674
rect 113100 73616 153106 73672
rect 153162 73616 153167 73672
rect 113100 73614 153167 73616
rect 113100 73612 113106 73614
rect 153101 73611 153167 73614
rect 161790 73612 161796 73676
rect 161860 73674 161866 73676
rect 194726 73674 194732 73676
rect 161860 73614 194732 73674
rect 161860 73612 161866 73614
rect 194726 73612 194732 73614
rect 194796 73612 194802 73676
rect 118374 73206 118802 73266
rect 116710 73068 116716 73132
rect 116780 73130 116786 73132
rect 118374 73130 118434 73206
rect 116780 73070 118434 73130
rect 118509 73132 118575 73133
rect 118509 73128 118556 73132
rect 118620 73130 118626 73132
rect 118742 73130 118802 73206
rect 156597 73132 156663 73133
rect 151118 73130 151124 73132
rect 118509 73072 118514 73128
rect 116780 73068 116786 73070
rect 118509 73068 118556 73072
rect 118620 73070 118666 73130
rect 118742 73070 151124 73130
rect 118620 73068 118626 73070
rect 151118 73068 151124 73070
rect 151188 73068 151194 73132
rect 156597 73128 156644 73132
rect 156708 73130 156714 73132
rect 170949 73130 171015 73133
rect 197302 73130 197308 73132
rect 156597 73072 156602 73128
rect 156597 73068 156644 73072
rect 156708 73070 156754 73130
rect 170949 73128 197308 73130
rect 170949 73072 170954 73128
rect 171010 73072 197308 73128
rect 170949 73070 197308 73072
rect 156708 73068 156714 73070
rect 118509 73067 118575 73068
rect 156597 73067 156663 73068
rect 170949 73067 171015 73070
rect 197302 73068 197308 73070
rect 197372 73068 197378 73132
rect 111006 72932 111012 72996
rect 111076 72994 111082 72996
rect 150433 72994 150499 72997
rect 111076 72992 150499 72994
rect 111076 72936 150438 72992
rect 150494 72936 150499 72992
rect 111076 72934 150499 72936
rect 111076 72932 111082 72934
rect 150433 72931 150499 72934
rect 173893 72994 173959 72997
rect 217041 72994 217107 72997
rect 173893 72992 217107 72994
rect 173893 72936 173898 72992
rect 173954 72936 217046 72992
rect 217102 72936 217107 72992
rect 173893 72934 217107 72936
rect 173893 72931 173959 72934
rect 217041 72931 217107 72934
rect 110873 72858 110939 72861
rect 142654 72858 142660 72860
rect 110873 72856 142660 72858
rect 110873 72800 110878 72856
rect 110934 72800 142660 72856
rect 110873 72798 142660 72800
rect 110873 72795 110939 72798
rect 142654 72796 142660 72798
rect 142724 72858 142730 72860
rect 165245 72858 165311 72861
rect 201534 72858 201540 72860
rect 142724 72798 147690 72858
rect 142724 72796 142730 72798
rect 104157 72722 104223 72725
rect 131021 72722 131087 72725
rect 104157 72720 131087 72722
rect 104157 72664 104162 72720
rect 104218 72664 131026 72720
rect 131082 72664 131087 72720
rect 104157 72662 131087 72664
rect 104157 72659 104223 72662
rect 131021 72659 131087 72662
rect 113582 72524 113588 72588
rect 113652 72586 113658 72588
rect 143809 72586 143875 72589
rect 113652 72584 143875 72586
rect 113652 72528 143814 72584
rect 143870 72528 143875 72584
rect 113652 72526 143875 72528
rect 113652 72524 113658 72526
rect 143809 72523 143875 72526
rect 115790 72388 115796 72452
rect 115860 72450 115866 72452
rect 145557 72450 145623 72453
rect 115860 72448 145623 72450
rect 115860 72392 145562 72448
rect 145618 72392 145623 72448
rect 115860 72390 145623 72392
rect 115860 72388 115866 72390
rect 145557 72387 145623 72390
rect -960 72178 480 72268
rect 113950 72252 113956 72316
rect 114020 72314 114026 72316
rect 139342 72314 139348 72316
rect 114020 72254 139348 72314
rect 114020 72252 114026 72254
rect 139342 72252 139348 72254
rect 139412 72252 139418 72316
rect 147630 72314 147690 72798
rect 165245 72856 201540 72858
rect 165245 72800 165250 72856
rect 165306 72800 201540 72856
rect 165245 72798 201540 72800
rect 165245 72795 165311 72798
rect 201534 72796 201540 72798
rect 201604 72796 201610 72860
rect 580257 72858 580323 72861
rect 583520 72858 584960 72948
rect 580257 72856 584960 72858
rect 580257 72800 580262 72856
rect 580318 72800 584960 72856
rect 580257 72798 584960 72800
rect 580257 72795 580323 72798
rect 158478 72660 158484 72724
rect 158548 72722 158554 72724
rect 192569 72722 192635 72725
rect 158548 72720 192635 72722
rect 158548 72664 192574 72720
rect 192630 72664 192635 72720
rect 583520 72708 584960 72798
rect 158548 72662 192635 72664
rect 158548 72660 158554 72662
rect 192569 72659 192635 72662
rect 164550 72524 164556 72588
rect 164620 72586 164626 72588
rect 198825 72586 198891 72589
rect 164620 72584 198891 72586
rect 164620 72528 198830 72584
rect 198886 72528 198891 72584
rect 164620 72526 198891 72528
rect 164620 72524 164626 72526
rect 198825 72523 198891 72526
rect 169661 72450 169727 72453
rect 191966 72450 191972 72452
rect 169661 72448 191972 72450
rect 169661 72392 169666 72448
rect 169722 72392 191972 72448
rect 169661 72390 191972 72392
rect 169661 72387 169727 72390
rect 191966 72388 191972 72390
rect 192036 72388 192042 72452
rect 580717 72314 580783 72317
rect 147630 72312 580783 72314
rect 147630 72256 580722 72312
rect 580778 72256 580783 72312
rect 147630 72254 580783 72256
rect 580717 72251 580783 72254
rect 3141 72178 3207 72181
rect -960 72176 3207 72178
rect -960 72120 3146 72176
rect 3202 72120 3207 72176
rect -960 72118 3207 72120
rect -960 72028 480 72118
rect 3141 72115 3207 72118
rect 123477 71770 123543 71773
rect 149646 71770 149652 71772
rect 123477 71768 149652 71770
rect 123477 71712 123482 71768
rect 123538 71712 149652 71768
rect 123477 71710 149652 71712
rect 123477 71707 123543 71710
rect 149646 71708 149652 71710
rect 149716 71708 149722 71772
rect 152457 71770 152523 71773
rect 152641 71770 152707 71773
rect 150758 71768 152707 71770
rect 150758 71712 152462 71768
rect 152518 71712 152646 71768
rect 152702 71712 152707 71768
rect 150758 71710 152707 71712
rect 118141 71634 118207 71637
rect 150758 71634 150818 71710
rect 152457 71707 152523 71710
rect 152641 71707 152707 71710
rect 156505 71770 156571 71773
rect 156689 71770 156755 71773
rect 187182 71770 187188 71772
rect 156505 71768 187188 71770
rect 156505 71712 156510 71768
rect 156566 71712 156694 71768
rect 156750 71712 187188 71768
rect 156505 71710 187188 71712
rect 156505 71707 156571 71710
rect 156689 71707 156755 71710
rect 187182 71708 187188 71710
rect 187252 71708 187258 71772
rect 118141 71632 150818 71634
rect 118141 71576 118146 71632
rect 118202 71576 150818 71632
rect 118141 71574 150818 71576
rect 159725 71634 159791 71637
rect 193438 71634 193444 71636
rect 159725 71632 193444 71634
rect 159725 71576 159730 71632
rect 159786 71576 193444 71632
rect 159725 71574 193444 71576
rect 118141 71571 118207 71574
rect 159725 71571 159791 71574
rect 193438 71572 193444 71574
rect 193508 71572 193514 71636
rect 112662 71436 112668 71500
rect 112732 71498 112738 71500
rect 147029 71498 147095 71501
rect 112732 71496 147095 71498
rect 112732 71440 147034 71496
rect 147090 71440 147095 71496
rect 112732 71438 147095 71440
rect 112732 71436 112738 71438
rect 147029 71435 147095 71438
rect 167678 71436 167684 71500
rect 167748 71498 167754 71500
rect 201493 71498 201559 71501
rect 167748 71496 201559 71498
rect 167748 71440 201498 71496
rect 201554 71440 201559 71496
rect 167748 71438 201559 71440
rect 167748 71436 167754 71438
rect 201493 71435 201559 71438
rect 207105 71498 207171 71501
rect 207606 71498 207612 71500
rect 207105 71496 207612 71498
rect 207105 71440 207110 71496
rect 207166 71440 207612 71496
rect 207105 71438 207612 71440
rect 207105 71435 207171 71438
rect 207606 71436 207612 71438
rect 207676 71436 207682 71500
rect 102910 71300 102916 71364
rect 102980 71362 102986 71364
rect 136582 71362 136588 71364
rect 102980 71302 136588 71362
rect 102980 71300 102986 71302
rect 136582 71300 136588 71302
rect 136652 71300 136658 71364
rect 171542 71300 171548 71364
rect 171612 71362 171618 71364
rect 205582 71362 205588 71364
rect 171612 71302 205588 71362
rect 171612 71300 171618 71302
rect 205582 71300 205588 71302
rect 205652 71300 205658 71364
rect 116853 71226 116919 71229
rect 149278 71226 149284 71228
rect 116853 71224 149284 71226
rect 116853 71168 116858 71224
rect 116914 71168 149284 71224
rect 116853 71166 149284 71168
rect 116853 71163 116919 71166
rect 149278 71164 149284 71166
rect 149348 71164 149354 71228
rect 173065 71226 173131 71229
rect 205766 71226 205772 71228
rect 173065 71224 205772 71226
rect 173065 71168 173070 71224
rect 173126 71168 205772 71224
rect 173065 71166 205772 71168
rect 173065 71163 173131 71166
rect 205766 71164 205772 71166
rect 205836 71164 205842 71228
rect 98545 71090 98611 71093
rect 156505 71090 156571 71093
rect 98545 71088 156571 71090
rect 98545 71032 98550 71088
rect 98606 71032 156510 71088
rect 156566 71032 156571 71088
rect 98545 71030 156571 71032
rect 98545 71027 98611 71030
rect 156505 71027 156571 71030
rect 166165 71090 166231 71093
rect 188102 71090 188108 71092
rect 166165 71088 188108 71090
rect 166165 71032 166170 71088
rect 166226 71032 188108 71088
rect 166165 71030 188108 71032
rect 166165 71027 166231 71030
rect 188102 71028 188108 71030
rect 188172 71028 188178 71092
rect 105721 70954 105787 70957
rect 133086 70954 133092 70956
rect 105721 70952 133092 70954
rect 105721 70896 105726 70952
rect 105782 70896 133092 70952
rect 105721 70894 133092 70896
rect 105721 70891 105787 70894
rect 133086 70892 133092 70894
rect 133156 70892 133162 70956
rect 162894 70892 162900 70956
rect 162964 70954 162970 70956
rect 218237 70954 218303 70957
rect 162964 70952 218303 70954
rect 162964 70896 218242 70952
rect 218298 70896 218303 70952
rect 162964 70894 218303 70896
rect 162964 70892 162970 70894
rect 218237 70891 218303 70894
rect 142061 70412 142127 70413
rect 142061 70408 142108 70412
rect 142172 70410 142178 70412
rect 142061 70352 142066 70408
rect 142061 70348 142108 70352
rect 142172 70350 142218 70410
rect 142172 70348 142178 70350
rect 142061 70347 142127 70348
rect 122598 70212 122604 70276
rect 122668 70274 122674 70276
rect 135897 70274 135963 70277
rect 122668 70272 135963 70274
rect 122668 70216 135902 70272
rect 135958 70216 135963 70272
rect 122668 70214 135963 70216
rect 122668 70212 122674 70214
rect 135897 70211 135963 70214
rect 165838 70212 165844 70276
rect 165908 70274 165914 70276
rect 186957 70274 187023 70277
rect 165908 70272 187023 70274
rect 165908 70216 186962 70272
rect 187018 70216 187023 70272
rect 165908 70214 187023 70216
rect 165908 70212 165914 70214
rect 186957 70211 187023 70214
rect 201493 70274 201559 70277
rect 202086 70274 202092 70276
rect 201493 70272 202092 70274
rect 201493 70216 201498 70272
rect 201554 70216 202092 70272
rect 201493 70214 202092 70216
rect 201493 70211 201559 70214
rect 202086 70212 202092 70214
rect 202156 70212 202162 70276
rect 204253 70274 204319 70277
rect 205030 70274 205036 70276
rect 204253 70272 205036 70274
rect 204253 70216 204258 70272
rect 204314 70216 205036 70272
rect 204253 70214 205036 70216
rect 204253 70211 204319 70214
rect 205030 70212 205036 70214
rect 205100 70212 205106 70276
rect 113766 70076 113772 70140
rect 113836 70138 113842 70140
rect 152181 70138 152247 70141
rect 113836 70136 152247 70138
rect 113836 70080 152186 70136
rect 152242 70080 152247 70136
rect 113836 70078 152247 70080
rect 113836 70076 113842 70078
rect 152181 70075 152247 70078
rect 175038 70076 175044 70140
rect 175108 70138 175114 70140
rect 207054 70138 207060 70140
rect 175108 70078 207060 70138
rect 175108 70076 175114 70078
rect 207054 70076 207060 70078
rect 207124 70076 207130 70140
rect 104566 69940 104572 70004
rect 104636 70002 104642 70004
rect 141693 70002 141759 70005
rect 104636 70000 141759 70002
rect 104636 69944 141698 70000
rect 141754 69944 141759 70000
rect 104636 69942 141759 69944
rect 104636 69940 104642 69942
rect 141693 69939 141759 69942
rect 170622 69940 170628 70004
rect 170692 70002 170698 70004
rect 204345 70002 204411 70005
rect 170692 70000 204411 70002
rect 170692 69944 204350 70000
rect 204406 69944 204411 70000
rect 170692 69942 204411 69944
rect 170692 69940 170698 69942
rect 204345 69939 204411 69942
rect 205633 70002 205699 70005
rect 206134 70002 206140 70004
rect 205633 70000 206140 70002
rect 205633 69944 205638 70000
rect 205694 69944 206140 70000
rect 205633 69942 206140 69944
rect 205633 69939 205699 69942
rect 206134 69940 206140 69942
rect 206204 69940 206210 70004
rect 100109 69866 100175 69869
rect 135294 69866 135300 69868
rect 100109 69864 135300 69866
rect 100109 69808 100114 69864
rect 100170 69808 135300 69864
rect 100109 69806 135300 69808
rect 100109 69803 100175 69806
rect 135294 69804 135300 69806
rect 135364 69804 135370 69868
rect 154246 69804 154252 69868
rect 154316 69866 154322 69868
rect 187734 69866 187740 69868
rect 154316 69806 187740 69866
rect 154316 69804 154322 69806
rect 187734 69804 187740 69806
rect 187804 69804 187810 69868
rect 112846 69668 112852 69732
rect 112916 69730 112922 69732
rect 145046 69730 145052 69732
rect 112916 69670 145052 69730
rect 112916 69668 112922 69670
rect 145046 69668 145052 69670
rect 145116 69668 145122 69732
rect 171317 69730 171383 69733
rect 196566 69730 196572 69732
rect 171317 69728 196572 69730
rect 171317 69672 171322 69728
rect 171378 69672 196572 69728
rect 171317 69670 196572 69672
rect 171317 69667 171383 69670
rect 196566 69668 196572 69670
rect 196636 69668 196642 69732
rect 108798 69532 108804 69596
rect 108868 69594 108874 69596
rect 139894 69594 139900 69596
rect 108868 69534 139900 69594
rect 108868 69532 108874 69534
rect 139894 69532 139900 69534
rect 139964 69532 139970 69596
rect 158294 69532 158300 69596
rect 158364 69594 158370 69596
rect 216949 69594 217015 69597
rect 158364 69592 217015 69594
rect 158364 69536 216954 69592
rect 217010 69536 217015 69592
rect 158364 69534 217015 69536
rect 158364 69532 158370 69534
rect 216949 69531 217015 69534
rect 108614 69396 108620 69460
rect 108684 69458 108690 69460
rect 150617 69458 150683 69461
rect 108684 69456 150683 69458
rect 108684 69400 150622 69456
rect 150678 69400 150683 69456
rect 108684 69398 150683 69400
rect 108684 69396 108690 69398
rect 150617 69395 150683 69398
rect 153469 69458 153535 69461
rect 187918 69458 187924 69460
rect 153469 69456 187924 69458
rect 153469 69400 153474 69456
rect 153530 69400 187924 69456
rect 153469 69398 187924 69400
rect 153469 69395 153535 69398
rect 187918 69396 187924 69398
rect 187988 69396 187994 69460
rect 121310 68852 121316 68916
rect 121380 68914 121386 68916
rect 135805 68914 135871 68917
rect 121380 68912 135871 68914
rect 121380 68856 135810 68912
rect 135866 68856 135871 68912
rect 121380 68854 135871 68856
rect 121380 68852 121386 68854
rect 135805 68851 135871 68854
rect 159357 68914 159423 68917
rect 205817 68914 205883 68917
rect 159357 68912 205883 68914
rect 159357 68856 159362 68912
rect 159418 68856 205822 68912
rect 205878 68856 205883 68912
rect 159357 68854 205883 68856
rect 159357 68851 159423 68854
rect 205817 68851 205883 68854
rect 106958 68716 106964 68780
rect 107028 68778 107034 68780
rect 141601 68778 141667 68781
rect 107028 68776 141667 68778
rect 107028 68720 141606 68776
rect 141662 68720 141667 68776
rect 107028 68718 141667 68720
rect 107028 68716 107034 68718
rect 141601 68715 141667 68718
rect 171133 68778 171199 68781
rect 209865 68778 209931 68781
rect 171133 68776 209931 68778
rect 171133 68720 171138 68776
rect 171194 68720 209870 68776
rect 209926 68720 209931 68776
rect 171133 68718 209931 68720
rect 171133 68715 171199 68718
rect 209865 68715 209931 68718
rect 579981 68778 580047 68781
rect 583520 68778 584960 68868
rect 579981 68776 584960 68778
rect 579981 68720 579986 68776
rect 580042 68720 584960 68776
rect 579981 68718 584960 68720
rect 579981 68715 580047 68718
rect 107326 68580 107332 68644
rect 107396 68642 107402 68644
rect 141509 68642 141575 68645
rect 107396 68640 141575 68642
rect 107396 68584 141514 68640
rect 141570 68584 141575 68640
rect 107396 68582 141575 68584
rect 107396 68580 107402 68582
rect 141509 68579 141575 68582
rect 168649 68642 168715 68645
rect 203006 68642 203012 68644
rect 168649 68640 203012 68642
rect 168649 68584 168654 68640
rect 168710 68584 203012 68640
rect 168649 68582 203012 68584
rect 168649 68579 168715 68582
rect 203006 68580 203012 68582
rect 203076 68580 203082 68644
rect 583520 68628 584960 68718
rect 111558 68444 111564 68508
rect 111628 68506 111634 68508
rect 143574 68506 143580 68508
rect 111628 68446 143580 68506
rect 111628 68444 111634 68446
rect 143574 68444 143580 68446
rect 143644 68444 143650 68508
rect 176510 68444 176516 68508
rect 176580 68506 176586 68508
rect 209814 68506 209820 68508
rect 176580 68446 209820 68506
rect 176580 68444 176586 68446
rect 209814 68444 209820 68446
rect 209884 68444 209890 68508
rect 107101 68370 107167 68373
rect 142061 68370 142127 68373
rect 107101 68368 142127 68370
rect 107101 68312 107106 68368
rect 107162 68312 142066 68368
rect 142122 68312 142127 68368
rect 107101 68310 142127 68312
rect 107101 68307 107167 68310
rect 142061 68307 142127 68310
rect 165337 68370 165403 68373
rect 172053 68370 172119 68373
rect 165337 68368 172119 68370
rect 165337 68312 165342 68368
rect 165398 68312 172058 68368
rect 172114 68312 172119 68368
rect 165337 68310 172119 68312
rect 165337 68307 165403 68310
rect 172053 68307 172119 68310
rect 173525 68370 173591 68373
rect 204621 68370 204687 68373
rect 173525 68368 204687 68370
rect 173525 68312 173530 68368
rect 173586 68312 204626 68368
rect 204682 68312 204687 68368
rect 173525 68310 204687 68312
rect 173525 68307 173591 68310
rect 204621 68307 204687 68310
rect 176469 68234 176535 68237
rect 206093 68234 206159 68237
rect 176469 68232 206159 68234
rect -960 68098 480 68188
rect 176469 68176 176474 68232
rect 176530 68176 206098 68232
rect 206154 68176 206159 68232
rect 176469 68174 206159 68176
rect 176469 68171 176535 68174
rect 206093 68171 206159 68174
rect 3141 68098 3207 68101
rect -960 68096 3207 68098
rect -960 68040 3146 68096
rect 3202 68040 3207 68096
rect -960 68038 3207 68040
rect -960 67948 480 68038
rect 3141 68035 3207 68038
rect 97717 67554 97783 67557
rect 138841 67554 138907 67557
rect 97717 67552 138907 67554
rect 97717 67496 97722 67552
rect 97778 67496 138846 67552
rect 138902 67496 138907 67552
rect 97717 67494 138907 67496
rect 97717 67491 97783 67494
rect 138841 67491 138907 67494
rect 163129 67554 163195 67557
rect 187366 67554 187372 67556
rect 163129 67552 187372 67554
rect 163129 67496 163134 67552
rect 163190 67496 187372 67552
rect 163129 67494 187372 67496
rect 163129 67491 163195 67494
rect 187366 67492 187372 67494
rect 187436 67492 187442 67556
rect 103278 67356 103284 67420
rect 103348 67418 103354 67420
rect 138238 67418 138244 67420
rect 103348 67358 138244 67418
rect 103348 67356 103354 67358
rect 138238 67356 138244 67358
rect 138308 67356 138314 67420
rect 174629 67418 174695 67421
rect 198958 67418 198964 67420
rect 174629 67416 198964 67418
rect 174629 67360 174634 67416
rect 174690 67360 198964 67416
rect 174629 67358 198964 67360
rect 174629 67355 174695 67358
rect 198958 67356 198964 67358
rect 199028 67356 199034 67420
rect 98913 67282 98979 67285
rect 132677 67282 132743 67285
rect 98913 67280 132743 67282
rect 98913 67224 98918 67280
rect 98974 67224 132682 67280
rect 132738 67224 132743 67280
rect 98913 67222 132743 67224
rect 98913 67219 98979 67222
rect 132677 67219 132743 67222
rect 166574 67220 166580 67284
rect 166644 67282 166650 67284
rect 201033 67282 201099 67285
rect 166644 67280 201099 67282
rect 166644 67224 201038 67280
rect 201094 67224 201099 67280
rect 166644 67222 201099 67224
rect 166644 67220 166650 67222
rect 201033 67219 201099 67222
rect 106038 67084 106044 67148
rect 106108 67146 106114 67148
rect 135846 67146 135852 67148
rect 106108 67086 135852 67146
rect 106108 67084 106114 67086
rect 135846 67084 135852 67086
rect 135916 67084 135922 67148
rect 167862 67084 167868 67148
rect 167932 67146 167938 67148
rect 201585 67146 201651 67149
rect 167932 67144 201651 67146
rect 167932 67088 201590 67144
rect 201646 67088 201651 67144
rect 167932 67086 201651 67088
rect 167932 67084 167938 67086
rect 201585 67083 201651 67086
rect 122966 66948 122972 67012
rect 123036 67010 123042 67012
rect 139761 67010 139827 67013
rect 123036 67008 139827 67010
rect 123036 66952 139766 67008
rect 139822 66952 139827 67008
rect 123036 66950 139827 66952
rect 123036 66948 123042 66950
rect 139761 66947 139827 66950
rect 162710 66948 162716 67012
rect 162780 67010 162786 67012
rect 192201 67010 192267 67013
rect 162780 67008 192267 67010
rect 162780 66952 192206 67008
rect 192262 66952 192267 67008
rect 162780 66950 192267 66952
rect 162780 66948 162786 66950
rect 192201 66947 192267 66950
rect 200205 67010 200271 67013
rect 200614 67010 200620 67012
rect 200205 67008 200620 67010
rect 200205 66952 200210 67008
rect 200266 66952 200620 67008
rect 200205 66950 200620 66952
rect 200205 66947 200271 66950
rect 200614 66948 200620 66950
rect 200684 66948 200690 67012
rect 170990 66812 170996 66876
rect 171060 66874 171066 66876
rect 211153 66874 211219 66877
rect 171060 66872 211219 66874
rect 171060 66816 211158 66872
rect 211214 66816 211219 66872
rect 171060 66814 211219 66816
rect 171060 66812 171066 66814
rect 211153 66811 211219 66814
rect 157425 66738 157491 66741
rect 192150 66738 192156 66740
rect 157425 66736 192156 66738
rect 157425 66680 157430 66736
rect 157486 66680 192156 66736
rect 157425 66678 192156 66680
rect 157425 66675 157491 66678
rect 192150 66676 192156 66678
rect 192220 66676 192226 66740
rect 103094 66132 103100 66196
rect 103164 66194 103170 66196
rect 136909 66194 136975 66197
rect 103164 66192 136975 66194
rect 103164 66136 136914 66192
rect 136970 66136 136975 66192
rect 103164 66134 136975 66136
rect 103164 66132 103170 66134
rect 136909 66131 136975 66134
rect 161054 66132 161060 66196
rect 161124 66194 161130 66196
rect 188981 66194 189047 66197
rect 161124 66192 189047 66194
rect 161124 66136 188986 66192
rect 189042 66136 189047 66192
rect 161124 66134 189047 66136
rect 161124 66132 161130 66134
rect 188981 66131 189047 66134
rect 107510 65996 107516 66060
rect 107580 66058 107586 66060
rect 140957 66058 141023 66061
rect 107580 66056 141023 66058
rect 107580 66000 140962 66056
rect 141018 66000 141023 66056
rect 107580 65998 141023 66000
rect 107580 65996 107586 65998
rect 140957 65995 141023 65998
rect 160686 65996 160692 66060
rect 160756 66058 160762 66060
rect 218145 66058 218211 66061
rect 160756 66056 218211 66058
rect 160756 66000 218150 66056
rect 218206 66000 218211 66056
rect 160756 65998 218211 66000
rect 160756 65996 160762 65998
rect 218145 65995 218211 65998
rect 104750 65860 104756 65924
rect 104820 65922 104826 65924
rect 138054 65922 138060 65924
rect 104820 65862 138060 65922
rect 104820 65860 104826 65862
rect 138054 65860 138060 65862
rect 138124 65860 138130 65924
rect 158110 65860 158116 65924
rect 158180 65922 158186 65924
rect 215753 65922 215819 65925
rect 158180 65920 215819 65922
rect 158180 65864 215758 65920
rect 215814 65864 215819 65920
rect 158180 65862 215819 65864
rect 158180 65860 158186 65862
rect 215753 65859 215819 65862
rect 108246 65724 108252 65788
rect 108316 65786 108322 65788
rect 140865 65786 140931 65789
rect 108316 65784 140931 65786
rect 108316 65728 140870 65784
rect 140926 65728 140931 65784
rect 108316 65726 140931 65728
rect 108316 65724 108322 65726
rect 140865 65723 140931 65726
rect 161974 65724 161980 65788
rect 162044 65786 162050 65788
rect 216857 65786 216923 65789
rect 162044 65784 216923 65786
rect 162044 65728 216862 65784
rect 216918 65728 216923 65784
rect 162044 65726 216923 65728
rect 162044 65724 162050 65726
rect 216857 65723 216923 65726
rect 164918 65588 164924 65652
rect 164988 65650 164994 65652
rect 199469 65650 199535 65653
rect 164988 65648 199535 65650
rect 164988 65592 199474 65648
rect 199530 65592 199535 65648
rect 164988 65590 199535 65592
rect 164988 65588 164994 65590
rect 199469 65587 199535 65590
rect 158989 65514 159055 65517
rect 186078 65514 186084 65516
rect 158989 65512 186084 65514
rect 158989 65456 158994 65512
rect 159050 65456 186084 65512
rect 158989 65454 186084 65456
rect 158989 65451 159055 65454
rect 186078 65452 186084 65454
rect 186148 65452 186154 65516
rect 154430 65316 154436 65380
rect 154500 65378 154506 65380
rect 214833 65378 214899 65381
rect 154500 65376 214899 65378
rect 154500 65320 214838 65376
rect 214894 65320 214899 65376
rect 154500 65318 214899 65320
rect 154500 65316 154506 65318
rect 214833 65315 214899 65318
rect 97625 64834 97691 64837
rect 144126 64834 144132 64836
rect 97625 64832 144132 64834
rect 97625 64776 97630 64832
rect 97686 64776 144132 64832
rect 97625 64774 144132 64776
rect 97625 64771 97691 64774
rect 144126 64772 144132 64774
rect 144196 64772 144202 64836
rect 158805 64834 158871 64837
rect 193254 64834 193260 64836
rect 158805 64832 193260 64834
rect 158805 64776 158810 64832
rect 158866 64776 193260 64832
rect 158805 64774 193260 64776
rect 158805 64771 158871 64774
rect 193254 64772 193260 64774
rect 193324 64772 193330 64836
rect 116894 64636 116900 64700
rect 116964 64698 116970 64700
rect 151169 64698 151235 64701
rect 116964 64696 151235 64698
rect 116964 64640 151174 64696
rect 151230 64640 151235 64696
rect 116964 64638 151235 64640
rect 116964 64636 116970 64638
rect 151169 64635 151235 64638
rect 169150 64636 169156 64700
rect 169220 64698 169226 64700
rect 200757 64698 200823 64701
rect 169220 64696 200823 64698
rect 169220 64640 200762 64696
rect 200818 64640 200823 64696
rect 169220 64638 200823 64640
rect 169220 64636 169226 64638
rect 200757 64635 200823 64638
rect 103329 64562 103395 64565
rect 134793 64562 134859 64565
rect 103329 64560 134859 64562
rect 103329 64504 103334 64560
rect 103390 64504 134798 64560
rect 134854 64504 134859 64560
rect 103329 64502 134859 64504
rect 103329 64499 103395 64502
rect 134793 64499 134859 64502
rect 163446 64500 163452 64564
rect 163516 64562 163522 64564
rect 194542 64562 194548 64564
rect 163516 64502 194548 64562
rect 163516 64500 163522 64502
rect 194542 64500 194548 64502
rect 194612 64500 194618 64564
rect 583520 64548 584960 64788
rect 119654 64364 119660 64428
rect 119724 64426 119730 64428
rect 147806 64426 147812 64428
rect 119724 64366 147812 64426
rect 119724 64364 119730 64366
rect 147806 64364 147812 64366
rect 147876 64364 147882 64428
rect 122046 64228 122052 64292
rect 122116 64290 122122 64292
rect 147990 64290 147996 64292
rect 122116 64230 147996 64290
rect 122116 64228 122122 64230
rect 147990 64228 147996 64230
rect 148060 64228 148066 64292
rect -960 64018 480 64108
rect 3141 64018 3207 64021
rect -960 64016 3207 64018
rect -960 63960 3146 64016
rect 3202 63960 3207 64016
rect -960 63958 3207 63960
rect -960 63868 480 63958
rect 3141 63955 3207 63958
rect 134793 63882 134859 63885
rect 134926 63882 134932 63884
rect 134793 63880 134932 63882
rect 134793 63824 134798 63880
rect 134854 63824 134932 63880
rect 134793 63822 134932 63824
rect 134793 63819 134859 63822
rect 134926 63820 134932 63822
rect 134996 63820 135002 63884
rect 161238 63412 161244 63476
rect 161308 63474 161314 63476
rect 211337 63474 211403 63477
rect 161308 63472 211403 63474
rect 161308 63416 211342 63472
rect 211398 63416 211403 63472
rect 161308 63414 211403 63416
rect 161308 63412 161314 63414
rect 211337 63411 211403 63414
rect 166758 63276 166764 63340
rect 166828 63338 166834 63340
rect 214189 63338 214255 63341
rect 166828 63336 214255 63338
rect 166828 63280 214194 63336
rect 214250 63280 214255 63336
rect 166828 63278 214255 63280
rect 166828 63276 166834 63278
rect 214189 63275 214255 63278
rect 168046 63140 168052 63204
rect 168116 63202 168122 63204
rect 211245 63202 211311 63205
rect 168116 63200 211311 63202
rect 168116 63144 211250 63200
rect 211306 63144 211311 63200
rect 168116 63142 211311 63144
rect 168116 63140 168122 63142
rect 211245 63139 211311 63142
rect 134926 62052 134932 62116
rect 134996 62114 135002 62116
rect 580441 62114 580507 62117
rect 134996 62112 580507 62114
rect 134996 62056 580446 62112
rect 580502 62056 580507 62112
rect 134996 62054 580507 62056
rect 134996 62052 135002 62054
rect 580441 62051 580507 62054
rect 583520 60468 584960 60708
rect -960 59788 480 60028
rect -960 56538 480 56628
rect 3417 56538 3483 56541
rect -960 56536 3483 56538
rect -960 56480 3422 56536
rect 3478 56480 3483 56536
rect -960 56478 3483 56480
rect -960 56388 480 56478
rect 3417 56475 3483 56478
rect 583520 56388 584960 56628
rect -960 52458 480 52548
rect 3417 52458 3483 52461
rect -960 52456 3483 52458
rect -960 52400 3422 52456
rect 3478 52400 3483 52456
rect -960 52398 3483 52400
rect -960 52308 480 52398
rect 3417 52395 3483 52398
rect 583520 52308 584960 52548
rect -960 48378 480 48468
rect 3233 48378 3299 48381
rect -960 48376 3299 48378
rect -960 48320 3238 48376
rect 3294 48320 3299 48376
rect -960 48318 3299 48320
rect -960 48228 480 48318
rect 3233 48315 3299 48318
rect 580165 48378 580231 48381
rect 583520 48378 584960 48468
rect 580165 48376 584960 48378
rect 580165 48320 580170 48376
rect 580226 48320 584960 48376
rect 580165 48318 584960 48320
rect 580165 48315 580231 48318
rect 583520 48228 584960 48318
rect -960 44298 480 44388
rect 3509 44298 3575 44301
rect -960 44296 3575 44298
rect -960 44240 3514 44296
rect 3570 44240 3575 44296
rect -960 44238 3575 44240
rect -960 44148 480 44238
rect 3509 44235 3575 44238
rect 579981 44298 580047 44301
rect 583520 44298 584960 44388
rect 579981 44296 584960 44298
rect 579981 44240 579986 44296
rect 580042 44240 584960 44296
rect 579981 44238 584960 44240
rect 579981 44235 580047 44238
rect 583520 44148 584960 44238
rect 580165 40898 580231 40901
rect 583520 40898 584960 40988
rect 580165 40896 584960 40898
rect 580165 40840 580170 40896
rect 580226 40840 584960 40896
rect 580165 40838 584960 40840
rect 580165 40835 580231 40838
rect 583520 40748 584960 40838
rect -960 40218 480 40308
rect 3509 40218 3575 40221
rect -960 40216 3575 40218
rect -960 40160 3514 40216
rect 3570 40160 3575 40216
rect -960 40158 3575 40160
rect -960 40068 480 40158
rect 3509 40155 3575 40158
rect 580165 36818 580231 36821
rect 583520 36818 584960 36908
rect 580165 36816 584960 36818
rect 580165 36760 580170 36816
rect 580226 36760 584960 36816
rect 580165 36758 584960 36760
rect 580165 36755 580231 36758
rect 583520 36668 584960 36758
rect -960 36138 480 36228
rect 3141 36138 3207 36141
rect -960 36136 3207 36138
rect -960 36080 3146 36136
rect 3202 36080 3207 36136
rect -960 36078 3207 36080
rect -960 35988 480 36078
rect 3141 36075 3207 36078
rect 580165 32738 580231 32741
rect 583520 32738 584960 32828
rect 580165 32736 584960 32738
rect 580165 32680 580170 32736
rect 580226 32680 584960 32736
rect 580165 32678 584960 32680
rect 580165 32675 580231 32678
rect 583520 32588 584960 32678
rect -960 32058 480 32148
rect 3141 32058 3207 32061
rect -960 32056 3207 32058
rect -960 32000 3146 32056
rect 3202 32000 3207 32056
rect -960 31998 3207 32000
rect -960 31908 480 31998
rect 3141 31995 3207 31998
rect 583520 28508 584960 28748
rect -960 27978 480 28068
rect 3141 27978 3207 27981
rect -960 27976 3207 27978
rect -960 27920 3146 27976
rect 3202 27920 3207 27976
rect -960 27918 3207 27920
rect -960 27828 480 27918
rect 3141 27915 3207 27918
rect 580165 24578 580231 24581
rect 583520 24578 584960 24668
rect 580165 24576 584960 24578
rect 580165 24520 580170 24576
rect 580226 24520 584960 24576
rect 580165 24518 584960 24520
rect 580165 24515 580231 24518
rect 583520 24428 584960 24518
rect -960 23898 480 23988
rect 3049 23898 3115 23901
rect -960 23896 3115 23898
rect -960 23840 3054 23896
rect 3110 23840 3115 23896
rect -960 23838 3115 23840
rect -960 23748 480 23838
rect 3049 23835 3115 23838
rect 580165 20498 580231 20501
rect 583520 20498 584960 20588
rect 580165 20496 584960 20498
rect 580165 20440 580170 20496
rect 580226 20440 584960 20496
rect 580165 20438 584960 20440
rect 580165 20435 580231 20438
rect 583520 20348 584960 20438
rect -960 19818 480 19908
rect 3509 19818 3575 19821
rect -960 19816 3575 19818
rect -960 19760 3514 19816
rect 3570 19760 3575 19816
rect -960 19758 3575 19760
rect -960 19668 480 19758
rect 3509 19755 3575 19758
rect 580165 16418 580231 16421
rect 583520 16418 584960 16508
rect 580165 16416 584960 16418
rect 580165 16360 580170 16416
rect 580226 16360 584960 16416
rect 580165 16358 584960 16360
rect 580165 16355 580231 16358
rect 583520 16268 584960 16358
rect -960 15738 480 15828
rect 3509 15738 3575 15741
rect -960 15736 3575 15738
rect -960 15680 3514 15736
rect 3570 15680 3575 15736
rect -960 15678 3575 15680
rect -960 15588 480 15678
rect 3509 15675 3575 15678
rect 580165 12338 580231 12341
rect 583520 12338 584960 12428
rect 580165 12336 584960 12338
rect 580165 12280 580170 12336
rect 580226 12280 584960 12336
rect 580165 12278 584960 12280
rect 580165 12275 580231 12278
rect 583520 12188 584960 12278
rect -960 11658 480 11748
rect 3049 11658 3115 11661
rect -960 11656 3115 11658
rect -960 11600 3054 11656
rect 3110 11600 3115 11656
rect -960 11598 3115 11600
rect -960 11508 480 11598
rect 3049 11595 3115 11598
rect 580165 8258 580231 8261
rect 583520 8258 584960 8348
rect 580165 8256 584960 8258
rect 580165 8200 580170 8256
rect 580226 8200 584960 8256
rect 580165 8198 584960 8200
rect 580165 8195 580231 8198
rect 583520 8108 584960 8198
rect -960 7578 480 7668
rect 2957 7578 3023 7581
rect -960 7576 3023 7578
rect -960 7520 2962 7576
rect 3018 7520 3023 7576
rect -960 7518 3023 7520
rect -960 7428 480 7518
rect 2957 7515 3023 7518
rect 580165 4178 580231 4181
rect 583520 4178 584960 4268
rect 580165 4176 584960 4178
rect 580165 4120 580170 4176
rect 580226 4120 584960 4176
rect 580165 4118 584960 4120
rect 580165 4115 580231 4118
rect 583520 4028 584960 4118
rect -960 3498 480 3588
rect 3141 3498 3207 3501
rect -960 3496 3207 3498
rect -960 3440 3146 3496
rect 3202 3440 3207 3496
rect -960 3438 3207 3440
rect -960 3348 480 3438
rect 3141 3435 3207 3438
rect 578877 98 578943 101
rect 583520 98 584960 188
rect 578877 96 584960 98
rect 578877 40 578882 96
rect 578938 40 584960 96
rect 578877 38 584960 40
rect 578877 35 578943 38
rect 583520 -52 584960 38
<< via3 >>
rect 196020 269724 196084 269788
rect 194548 268364 194612 268428
rect 111748 265508 111812 265572
rect 118556 263876 118620 263940
rect 116900 263740 116964 263804
rect 196204 263604 196268 263668
rect 191788 262924 191852 262988
rect 111748 262788 111812 262852
rect 112852 262788 112916 262852
rect 193260 262788 193324 262852
rect 194548 262788 194612 262852
rect 196020 262516 196084 262580
rect 197492 262380 197556 262444
rect 121500 262304 121564 262308
rect 121500 262248 121550 262304
rect 121550 262248 121564 262304
rect 121500 262244 121564 262248
rect 121316 260068 121380 260132
rect 122604 259992 122668 259996
rect 122604 259936 122618 259992
rect 122618 259936 122668 259992
rect 122604 259932 122668 259936
rect 187188 259932 187252 259996
rect 111564 259660 111628 259724
rect 111380 259524 111444 259588
rect 187004 259312 187068 259316
rect 187004 259256 187018 259312
rect 187018 259256 187068 259312
rect 187004 259252 187068 259256
rect 188292 245652 188356 245716
rect 122052 237356 122116 237420
rect 186820 233276 186884 233340
rect 121500 218044 121564 218108
rect 188476 218044 188540 218108
rect 122236 216684 122300 216748
rect 122420 212604 122484 212668
rect 138612 201452 138676 201516
rect 160324 201452 160388 201516
rect 181484 201724 181548 201788
rect 184980 201452 185044 201516
rect 207060 201044 207124 201108
rect 154252 200908 154316 200972
rect 180196 200908 180260 200972
rect 186820 200908 186884 200972
rect 205036 200908 205100 200972
rect 122236 200772 122300 200836
rect 146524 200772 146588 200836
rect 188292 200772 188356 200836
rect 210924 200772 210988 200836
rect 137876 200636 137940 200700
rect 211108 200636 211172 200700
rect 173572 200500 173636 200564
rect 205036 200500 205100 200564
rect 122052 200364 122116 200428
rect 140452 200228 140516 200292
rect 170628 200364 170692 200428
rect 158116 200228 158180 200292
rect 160876 200228 160940 200292
rect 169524 200228 169588 200292
rect 207060 200364 207124 200428
rect 211108 200228 211172 200292
rect 133644 199820 133708 199884
rect 133828 199858 133832 199884
rect 133832 199858 133888 199884
rect 133888 199858 133892 199884
rect 133828 199820 133892 199858
rect 134196 199880 134260 199884
rect 134196 199824 134200 199880
rect 134200 199824 134256 199880
rect 134256 199824 134260 199880
rect 134196 199820 134260 199824
rect 135116 199858 135120 199884
rect 135120 199858 135176 199884
rect 135176 199858 135180 199884
rect 135116 199820 135180 199858
rect 136220 199820 136284 199884
rect 136404 199684 136468 199748
rect 135852 199548 135916 199612
rect 138428 199880 138492 199884
rect 138428 199824 138432 199880
rect 138432 199824 138488 199880
rect 138488 199824 138492 199880
rect 138428 199820 138492 199824
rect 138796 199820 138860 199884
rect 139348 199880 139412 199884
rect 139348 199824 139352 199880
rect 139352 199824 139408 199880
rect 139408 199824 139412 199880
rect 139348 199820 139412 199824
rect 140084 199880 140148 199884
rect 140084 199824 140088 199880
rect 140088 199824 140144 199880
rect 140144 199824 140148 199880
rect 140084 199820 140148 199824
rect 140268 199880 140332 199884
rect 140268 199824 140272 199880
rect 140272 199824 140328 199880
rect 140328 199824 140332 199880
rect 140268 199820 140332 199824
rect 141004 199820 141068 199884
rect 142476 199880 142540 199884
rect 142476 199824 142480 199880
rect 142480 199824 142536 199880
rect 142536 199824 142540 199880
rect 142476 199820 142540 199824
rect 144684 199820 144748 199884
rect 145236 199820 145300 199884
rect 146524 199820 146588 199884
rect 138244 199684 138308 199748
rect 138612 199684 138676 199748
rect 139716 199684 139780 199748
rect 141372 199684 141436 199748
rect 143028 199684 143092 199748
rect 143948 199684 144012 199748
rect 147444 199820 147508 199884
rect 147996 199820 148060 199884
rect 148180 199684 148244 199748
rect 143212 199548 143276 199612
rect 143580 199548 143644 199612
rect 146892 199548 146956 199612
rect 152596 200092 152660 200156
rect 149468 199880 149532 199884
rect 149468 199824 149472 199880
rect 149472 199824 149528 199880
rect 149528 199824 149532 199880
rect 149468 199820 149532 199824
rect 150020 199820 150084 199884
rect 150572 199820 150636 199884
rect 151124 199820 151188 199884
rect 151860 199744 151924 199748
rect 151860 199688 151910 199744
rect 151910 199688 151924 199744
rect 151860 199684 151924 199688
rect 152228 199684 152292 199748
rect 152964 199858 152968 199884
rect 152968 199858 153024 199884
rect 153024 199858 153028 199884
rect 152964 199820 153028 199858
rect 153884 199820 153948 199884
rect 154068 199820 154132 199884
rect 157012 199880 157076 199884
rect 157012 199824 157016 199880
rect 157016 199824 157072 199880
rect 157072 199824 157076 199880
rect 157012 199820 157076 199824
rect 157380 199820 157444 199884
rect 163452 200092 163516 200156
rect 158300 199858 158304 199884
rect 158304 199858 158360 199884
rect 158360 199858 158364 199884
rect 158300 199820 158364 199858
rect 151308 199548 151372 199612
rect 156828 199744 156892 199748
rect 156828 199688 156842 199744
rect 156842 199688 156892 199744
rect 156828 199684 156892 199688
rect 158116 199684 158180 199748
rect 152964 199608 153028 199612
rect 152964 199552 152978 199608
rect 152978 199552 153028 199608
rect 152964 199548 153028 199552
rect 153332 199608 153396 199612
rect 153332 199552 153382 199608
rect 153382 199552 153396 199608
rect 153332 199548 153396 199552
rect 154252 199548 154316 199612
rect 156644 199548 156708 199612
rect 159404 199820 159468 199884
rect 160324 199820 160388 199884
rect 159588 199684 159652 199748
rect 161980 199820 162044 199884
rect 163268 199956 163332 200020
rect 164004 199880 164068 199884
rect 164004 199824 164008 199880
rect 164008 199824 164064 199880
rect 164064 199824 164068 199880
rect 164004 199820 164068 199824
rect 164556 199820 164620 199884
rect 166580 199956 166644 200020
rect 166396 199820 166460 199884
rect 162532 199684 162596 199748
rect 166028 199684 166092 199748
rect 166212 199684 166276 199748
rect 167316 199858 167320 199884
rect 167320 199858 167376 199884
rect 167376 199858 167380 199884
rect 167316 199820 167380 199858
rect 168604 199880 168668 199884
rect 168604 199824 168608 199880
rect 168608 199824 168664 199880
rect 168664 199824 168668 199880
rect 168604 199820 168668 199824
rect 168972 199820 169036 199884
rect 169340 199684 169404 199748
rect 170996 200092 171060 200156
rect 173204 199956 173268 200020
rect 170628 199858 170632 199884
rect 170632 199858 170688 199884
rect 170688 199858 170692 199884
rect 170628 199820 170692 199858
rect 171364 199820 171428 199884
rect 172284 199820 172348 199884
rect 174308 199858 174312 199884
rect 174312 199858 174368 199884
rect 174368 199858 174372 199884
rect 174308 199820 174372 199858
rect 174676 199858 174680 199884
rect 174680 199858 174736 199884
rect 174736 199858 174740 199884
rect 174676 199820 174740 199858
rect 209820 200092 209884 200156
rect 210924 200092 210988 200156
rect 180196 199956 180260 200020
rect 176332 199820 176396 199884
rect 188476 199684 188540 199748
rect 160876 199548 160940 199612
rect 164740 199548 164804 199612
rect 165108 199548 165172 199612
rect 169156 199548 169220 199612
rect 169524 199548 169588 199612
rect 170812 199608 170876 199612
rect 170812 199552 170862 199608
rect 170862 199552 170876 199608
rect 170812 199548 170876 199552
rect 205588 199548 205652 199612
rect 107516 199412 107580 199476
rect 122420 199412 122484 199476
rect 175412 199412 175476 199476
rect 176332 199412 176396 199476
rect 161980 199276 162044 199340
rect 163268 199276 163332 199340
rect 168420 199276 168484 199340
rect 139716 199140 139780 199204
rect 140084 199200 140148 199204
rect 140084 199144 140098 199200
rect 140098 199144 140148 199200
rect 140084 199140 140148 199144
rect 140452 199140 140516 199204
rect 153700 199140 153764 199204
rect 184980 199140 185044 199204
rect 143396 199004 143460 199068
rect 150572 199004 150636 199068
rect 151492 199004 151556 199068
rect 151676 199064 151740 199068
rect 151676 199008 151690 199064
rect 151690 199008 151740 199064
rect 151676 199004 151740 199008
rect 151124 198868 151188 198932
rect 151308 198868 151372 198932
rect 152044 198868 152108 198932
rect 153884 198868 153948 198932
rect 158300 198868 158364 198932
rect 167868 198868 167932 198932
rect 173572 198868 173636 198932
rect 205588 198868 205652 198932
rect 206140 198868 206204 198932
rect 107516 198732 107580 198796
rect 164740 198732 164804 198796
rect 138796 198596 138860 198660
rect 162716 198596 162780 198660
rect 173388 198596 173452 198660
rect 173756 198656 173820 198660
rect 173756 198600 173770 198656
rect 173770 198600 173820 198656
rect 173756 198596 173820 198600
rect 174676 198656 174740 198660
rect 174676 198600 174690 198656
rect 174690 198600 174740 198656
rect 174676 198596 174740 198600
rect 140268 198460 140332 198524
rect 142292 198520 142356 198524
rect 142292 198464 142306 198520
rect 142306 198464 142356 198520
rect 142292 198460 142356 198464
rect 144500 198460 144564 198524
rect 147076 198324 147140 198388
rect 165476 198324 165540 198388
rect 138980 198188 139044 198252
rect 141372 198188 141436 198252
rect 159588 198188 159652 198252
rect 134380 197780 134444 197844
rect 147996 197916 148060 197980
rect 148916 197976 148980 197980
rect 148916 197920 148966 197976
rect 148966 197920 148980 197976
rect 148916 197916 148980 197920
rect 163636 197916 163700 197980
rect 185348 197916 185412 197980
rect 141004 197780 141068 197844
rect 157012 197780 157076 197844
rect 164004 197780 164068 197844
rect 168236 197644 168300 197708
rect 145236 197508 145300 197572
rect 169708 197508 169772 197572
rect 171364 197508 171428 197572
rect 142476 197372 142540 197436
rect 151124 197372 151188 197436
rect 170812 197432 170876 197436
rect 170812 197376 170826 197432
rect 170826 197376 170876 197432
rect 170812 197372 170876 197376
rect 176516 197372 176580 197436
rect 132540 197100 132604 197164
rect 133644 197100 133708 197164
rect 141004 197100 141068 197164
rect 144132 197100 144196 197164
rect 147444 197100 147508 197164
rect 164004 196964 164068 197028
rect 173388 197024 173452 197028
rect 173388 196968 173402 197024
rect 173402 196968 173452 197024
rect 173388 196964 173452 196968
rect 210372 196964 210436 197028
rect 210924 196964 210988 197028
rect 122236 196692 122300 196756
rect 138244 196752 138308 196756
rect 138244 196696 138258 196752
rect 138258 196696 138308 196752
rect 138244 196692 138308 196696
rect 139900 196692 139964 196756
rect 143212 196692 143276 196756
rect 149100 196752 149164 196756
rect 149100 196696 149150 196752
rect 149150 196696 149164 196752
rect 149100 196692 149164 196696
rect 151860 196692 151924 196756
rect 157196 196692 157260 196756
rect 161244 196752 161308 196756
rect 161244 196696 161258 196752
rect 161258 196696 161308 196752
rect 161244 196692 161308 196696
rect 163820 196692 163884 196756
rect 164372 196692 164436 196756
rect 170996 196692 171060 196756
rect 205588 196692 205652 196756
rect 210924 196692 210988 196756
rect 117084 196556 117148 196620
rect 149468 196556 149532 196620
rect 190500 196556 190564 196620
rect 133828 196420 133892 196484
rect 137876 196420 137940 196484
rect 138796 196420 138860 196484
rect 157380 196420 157444 196484
rect 171732 196420 171796 196484
rect 135116 196284 135180 196348
rect 167316 196284 167380 196348
rect 137324 196208 137388 196212
rect 137324 196152 137374 196208
rect 137374 196152 137388 196208
rect 137324 196148 137388 196152
rect 137876 196148 137940 196212
rect 154068 196148 154132 196212
rect 139348 196012 139412 196076
rect 152596 196072 152660 196076
rect 152596 196016 152646 196072
rect 152646 196016 152660 196072
rect 152596 196012 152660 196016
rect 153884 196012 153948 196076
rect 154252 196012 154316 196076
rect 156644 196012 156708 196076
rect 174676 196012 174740 196076
rect 122604 195876 122668 195940
rect 136036 195876 136100 195940
rect 136404 195936 136468 195940
rect 136404 195880 136454 195936
rect 136454 195880 136468 195936
rect 136404 195876 136468 195880
rect 137140 195876 137204 195940
rect 138428 195936 138492 195940
rect 138428 195880 138442 195936
rect 138442 195880 138492 195936
rect 138428 195876 138492 195880
rect 138612 195876 138676 195940
rect 143948 195876 144012 195940
rect 174860 195740 174924 195804
rect 124076 195604 124140 195668
rect 164556 195392 164620 195396
rect 164556 195336 164570 195392
rect 164570 195336 164620 195392
rect 164556 195332 164620 195336
rect 165476 195332 165540 195396
rect 168604 195196 168668 195260
rect 143028 195120 143092 195124
rect 143028 195064 143042 195120
rect 143042 195064 143092 195120
rect 143028 195060 143092 195064
rect 214052 195060 214116 195124
rect 121316 194576 121380 194580
rect 121316 194520 121366 194576
rect 121366 194520 121380 194576
rect 121316 194516 121380 194520
rect 108804 194108 108868 194172
rect 142292 194108 142356 194172
rect 99236 193972 99300 194036
rect 197308 193972 197372 194036
rect 119660 193836 119724 193900
rect 198780 193836 198844 193900
rect 146708 193760 146772 193764
rect 146708 193704 146722 193760
rect 146722 193704 146772 193760
rect 146708 193700 146772 193704
rect 154068 193760 154132 193764
rect 154068 193704 154118 193760
rect 154118 193704 154132 193760
rect 154068 193700 154132 193704
rect 134196 193292 134260 193356
rect 175228 193156 175292 193220
rect 173020 193020 173084 193084
rect 205772 193020 205836 193084
rect 119660 192884 119724 192948
rect 149100 192884 149164 192948
rect 164372 192884 164436 192948
rect 168420 192748 168484 192812
rect 166396 192476 166460 192540
rect 200620 192476 200684 192540
rect 153148 191660 153212 191724
rect 167868 191524 167932 191588
rect 202092 191524 202156 191588
rect 166580 191252 166644 191316
rect 122604 191116 122668 191180
rect 156828 191116 156892 191180
rect 114140 190980 114204 191044
rect 161244 190980 161308 191044
rect 166028 190844 166092 190908
rect 189028 190708 189092 190772
rect 163820 190572 163884 190636
rect 197308 190572 197372 190636
rect 113036 190436 113100 190500
rect 137324 190360 137388 190364
rect 137324 190304 137338 190360
rect 137338 190304 137388 190360
rect 137324 190300 137388 190304
rect 148180 190300 148244 190364
rect 175412 190164 175476 190228
rect 163452 190028 163516 190092
rect 191972 190028 192036 190092
rect 193076 190028 193140 190092
rect 187740 189892 187804 189956
rect 119660 189756 119724 189820
rect 172284 189756 172348 189820
rect 118372 189620 118436 189684
rect 187740 189620 187804 189684
rect 193076 189620 193140 189684
rect 148180 189076 148244 189140
rect 151124 189076 151188 189140
rect 163636 189136 163700 189140
rect 163636 189080 163650 189136
rect 163650 189080 163700 189136
rect 163636 189076 163700 189080
rect 175412 189136 175476 189140
rect 175412 189080 175462 189136
rect 175462 189080 175476 189136
rect 175412 189076 175476 189080
rect 144500 188940 144564 189004
rect 143396 188728 143460 188732
rect 143396 188672 143446 188728
rect 143446 188672 143460 188728
rect 143396 188668 143460 188672
rect 122420 188532 122484 188596
rect 132540 188396 132604 188460
rect 176516 188532 176580 188596
rect 162532 188396 162596 188460
rect 201540 188396 201604 188460
rect 143580 188260 143644 188324
rect 151492 188260 151556 188324
rect 169708 187580 169772 187644
rect 147076 187444 147140 187508
rect 122972 187308 123036 187372
rect 174676 187308 174740 187372
rect 207612 187308 207676 187372
rect 113956 187172 114020 187236
rect 174860 187172 174924 187236
rect 108436 187036 108500 187100
rect 168236 187036 168300 187100
rect 112484 186900 112548 186964
rect 147076 186900 147140 186964
rect 187924 186900 187988 186964
rect 169340 186764 169404 186828
rect 144132 186220 144196 186284
rect 146892 186220 146956 186284
rect 175228 186084 175292 186148
rect 169156 185948 169220 186012
rect 173756 185812 173820 185876
rect 174492 185676 174556 185740
rect 112668 185540 112732 185604
rect 146892 185540 146956 185604
rect 148916 185540 148980 185604
rect 189212 185540 189276 185604
rect 162716 184452 162780 184516
rect 164004 184316 164068 184380
rect 168972 184180 169036 184244
rect 203564 184180 203628 184244
rect 138980 183560 139044 183564
rect 138980 183504 139030 183560
rect 139030 183504 139044 183560
rect 138980 183500 139044 183504
rect 107148 182820 107212 182884
rect 139900 182820 139964 182884
rect 144684 183364 144748 183428
rect 159036 183228 159100 183292
rect 154068 183092 154132 183156
rect 185716 182956 185780 183020
rect 154252 182820 154316 182884
rect 186084 182820 186148 182884
rect 157196 182548 157260 182612
rect 108620 182140 108684 182204
rect 150020 182004 150084 182068
rect 151676 181324 151740 181388
rect 100524 180916 100588 180980
rect 104572 180780 104636 180844
rect 138796 180780 138860 180844
rect 137876 180644 137940 180708
rect 138796 180372 138860 180436
rect 104756 180100 104820 180164
rect 138612 180100 138676 180164
rect 107332 179964 107396 180028
rect 106044 179692 106108 179756
rect 103284 179556 103348 179620
rect 99052 179420 99116 179484
rect 136220 179420 136284 179484
rect 137876 179420 137940 179484
rect 166212 178876 166276 178940
rect 171732 178740 171796 178804
rect 203012 178740 203076 178804
rect 165108 178604 165172 178668
rect 141004 177924 141068 177988
rect 136036 177788 136100 177852
rect 122236 176564 122300 176628
rect 121132 176428 121196 176492
rect 102916 176292 102980 176356
rect 137140 176292 137204 176356
rect 103100 176156 103164 176220
rect 124812 176020 124876 176084
rect 121316 175884 121380 175948
rect 135852 175884 135916 175948
rect 100340 148548 100404 148612
rect 111012 148412 111076 148476
rect 106964 148276 107028 148340
rect 198964 146916 199028 146980
rect 111564 145964 111628 146028
rect 197492 145964 197556 146028
rect 111380 145828 111444 145892
rect 112852 145692 112916 145756
rect 196204 145692 196268 145756
rect 111564 144332 111628 144396
rect 196572 144332 196636 144396
rect 116532 144196 116596 144260
rect 161980 144196 162044 144260
rect 113772 144060 113836 144124
rect 192156 144060 192220 144124
rect 187188 143380 187252 143444
rect 196020 143244 196084 143308
rect 187004 143108 187068 143172
rect 116900 142972 116964 143036
rect 118556 142836 118620 142900
rect 193260 142836 193324 142900
rect 191788 142700 191852 142764
rect 112852 141884 112916 141948
rect 118556 141612 118620 141676
rect 193444 141612 193508 141676
rect 118188 141476 118252 141540
rect 196388 141476 196452 141540
rect 116716 141340 116780 141404
rect 181484 141340 181548 141404
rect 194548 141340 194612 141404
rect 120948 140660 121012 140724
rect 115612 140524 115676 140588
rect 193628 140524 193692 140588
rect 113588 140388 113652 140452
rect 134380 140252 134444 140316
rect 194732 140252 194796 140316
rect 120580 140116 120644 140180
rect 187372 140116 187436 140180
rect 121868 139980 121932 140044
rect 188108 139980 188172 140044
rect 196204 139980 196268 140044
rect 115428 139844 115492 139908
rect 187556 139708 187620 139772
rect 116900 139436 116964 139500
rect 122052 139300 122116 139364
rect 123892 139300 123956 139364
rect 126100 139300 126164 139364
rect 136956 139300 137020 139364
rect 108252 138756 108316 138820
rect 136956 138756 137020 138820
rect 187188 139300 187252 139364
rect 187004 139164 187068 139228
rect 190684 138892 190748 138956
rect 193812 138756 193876 138820
rect 126100 138484 126164 138548
rect 185348 138212 185412 138276
rect 186268 138212 186332 138276
rect 115796 138136 115860 138140
rect 115796 138080 115846 138136
rect 115846 138080 115860 138136
rect 115796 138076 115860 138080
rect 122972 137940 123036 138004
rect 111196 137804 111260 137868
rect 124812 137804 124876 137868
rect 185716 137804 185780 137868
rect 193260 137804 193324 137868
rect 187188 137396 187252 137460
rect 187556 137260 187620 137324
rect 186820 136580 186884 136644
rect 186268 134404 186332 134468
rect 122052 132636 122116 132700
rect 122788 132636 122852 132700
rect 122052 132364 122116 132428
rect 122788 132364 122852 132428
rect 122052 122980 122116 123044
rect 122788 122980 122852 123044
rect 122788 122708 122852 122772
rect 122788 113188 122852 113252
rect 122788 113052 122852 113116
rect 122788 103532 122852 103596
rect 122788 103396 122852 103460
rect 122788 93876 122852 93940
rect 122788 93740 122852 93804
rect 120580 92516 120644 92580
rect 186084 91156 186148 91220
rect 122972 83404 123036 83468
rect 187188 82724 187252 82788
rect 186084 82180 186148 82244
rect 193812 82180 193876 82244
rect 135852 81908 135916 81972
rect 176700 81908 176764 81972
rect 137324 81772 137388 81836
rect 175044 81772 175108 81836
rect 111196 81636 111260 81700
rect 119660 81500 119724 81564
rect 184796 81636 184860 81700
rect 141372 81364 141436 81428
rect 196388 81364 196452 81428
rect 131436 81228 131500 81292
rect 166580 81228 166644 81292
rect 133276 81092 133340 81156
rect 174860 81092 174924 81156
rect 203564 81092 203628 81156
rect 135484 80956 135548 81020
rect 166948 80956 167012 81020
rect 112484 80820 112548 80884
rect 147444 80820 147508 80884
rect 154804 80820 154868 80884
rect 99052 80684 99116 80748
rect 134380 80684 134444 80748
rect 116532 80548 116596 80612
rect 131436 80004 131500 80068
rect 133276 79868 133340 79932
rect 177252 80548 177316 80612
rect 190684 80548 190748 80612
rect 154252 80140 154316 80204
rect 161060 80140 161124 80204
rect 169156 80140 169220 80204
rect 186820 80004 186884 80068
rect 134380 79928 134444 79932
rect 134380 79872 134384 79928
rect 134384 79872 134440 79928
rect 134440 79872 134444 79928
rect 134380 79868 134444 79872
rect 135116 79928 135180 79932
rect 135116 79872 135120 79928
rect 135120 79872 135176 79928
rect 135176 79872 135180 79928
rect 135116 79868 135180 79872
rect 135668 79868 135732 79932
rect 136404 79906 136408 79932
rect 136408 79906 136464 79932
rect 136464 79906 136468 79932
rect 136404 79868 136468 79906
rect 134932 79792 134996 79796
rect 134932 79736 134936 79792
rect 134936 79736 134992 79792
rect 134992 79736 134996 79792
rect 134932 79732 134996 79736
rect 135300 79792 135364 79796
rect 135300 79736 135304 79792
rect 135304 79736 135360 79792
rect 135360 79736 135364 79792
rect 135300 79732 135364 79736
rect 135852 79792 135916 79796
rect 135852 79736 135902 79792
rect 135902 79736 135916 79792
rect 135852 79732 135916 79736
rect 136220 79732 136284 79796
rect 137324 79906 137328 79932
rect 137328 79906 137384 79932
rect 137384 79906 137388 79932
rect 137324 79868 137388 79906
rect 138612 79906 138616 79932
rect 138616 79906 138672 79932
rect 138672 79906 138676 79932
rect 138612 79868 138676 79906
rect 140084 79928 140148 79932
rect 140084 79872 140088 79928
rect 140088 79872 140144 79928
rect 140144 79872 140148 79928
rect 139348 79792 139412 79796
rect 139348 79736 139362 79792
rect 139362 79736 139412 79792
rect 139348 79732 139412 79736
rect 138060 79460 138124 79524
rect 122420 79324 122484 79388
rect 135116 79052 135180 79116
rect 135484 79052 135548 79116
rect 136772 79052 136836 79116
rect 138612 79324 138676 79388
rect 140084 79868 140148 79872
rect 140268 79906 140272 79932
rect 140272 79906 140328 79932
rect 140328 79906 140332 79932
rect 140268 79868 140332 79906
rect 141188 79868 141252 79932
rect 140636 79732 140700 79796
rect 144500 79868 144564 79932
rect 141372 79656 141436 79660
rect 141372 79600 141422 79656
rect 141422 79600 141436 79656
rect 141372 79596 141436 79600
rect 143948 79596 144012 79660
rect 145052 79656 145116 79660
rect 145052 79600 145102 79656
rect 145102 79600 145116 79656
rect 145052 79596 145116 79600
rect 147444 79906 147448 79932
rect 147448 79906 147504 79932
rect 147504 79906 147508 79932
rect 147444 79868 147508 79906
rect 148548 79928 148612 79932
rect 148548 79872 148552 79928
rect 148552 79872 148608 79928
rect 148608 79872 148612 79928
rect 148548 79868 148612 79872
rect 149468 79906 149472 79932
rect 149472 79906 149528 79932
rect 149528 79906 149532 79932
rect 149468 79868 149532 79906
rect 150940 79868 151004 79932
rect 147812 79324 147876 79388
rect 151124 79732 151188 79796
rect 152596 79928 152660 79932
rect 152596 79872 152600 79928
rect 152600 79872 152656 79928
rect 152656 79872 152660 79928
rect 152596 79868 152660 79872
rect 152780 79868 152844 79932
rect 153700 79906 153704 79932
rect 153704 79906 153760 79932
rect 153760 79906 153764 79932
rect 153700 79868 153764 79906
rect 154068 79928 154132 79932
rect 154068 79872 154072 79928
rect 154072 79872 154128 79928
rect 154128 79872 154132 79928
rect 154068 79868 154132 79872
rect 154252 79732 154316 79796
rect 139348 79248 139412 79252
rect 139348 79192 139362 79248
rect 139362 79192 139412 79248
rect 139348 79188 139412 79192
rect 154804 79656 154868 79660
rect 154804 79600 154818 79656
rect 154818 79600 154868 79656
rect 154804 79596 154868 79600
rect 158484 79732 158548 79796
rect 158852 79792 158916 79796
rect 158852 79736 158856 79792
rect 158856 79736 158912 79792
rect 158912 79736 158916 79792
rect 158852 79732 158916 79736
rect 159588 79732 159652 79796
rect 160508 79868 160572 79932
rect 161796 79868 161860 79932
rect 162348 79868 162412 79932
rect 163452 79906 163456 79932
rect 163456 79906 163512 79932
rect 163512 79906 163516 79932
rect 163452 79868 163516 79906
rect 163636 79732 163700 79796
rect 164556 79732 164620 79796
rect 166764 79868 166828 79932
rect 167132 79868 167196 79932
rect 167868 79928 167932 79932
rect 167868 79872 167872 79928
rect 167872 79872 167928 79928
rect 167928 79872 167932 79928
rect 167868 79868 167932 79872
rect 168236 79928 168300 79932
rect 168236 79872 168240 79928
rect 168240 79872 168296 79928
rect 168296 79872 168300 79928
rect 168236 79868 168300 79872
rect 166948 79792 167012 79796
rect 166948 79736 166952 79792
rect 166952 79736 167008 79792
rect 167008 79736 167012 79792
rect 166948 79732 167012 79736
rect 166396 79596 166460 79660
rect 166580 79656 166644 79660
rect 167684 79732 167748 79796
rect 166580 79600 166594 79656
rect 166594 79600 166644 79656
rect 166580 79596 166644 79600
rect 168052 79596 168116 79660
rect 170076 79868 170140 79932
rect 172284 79906 172288 79932
rect 172288 79906 172344 79932
rect 172344 79906 172348 79932
rect 172284 79868 172348 79906
rect 170628 79732 170692 79796
rect 170812 79732 170876 79796
rect 171548 79792 171612 79796
rect 171548 79736 171598 79792
rect 171598 79736 171612 79792
rect 171548 79732 171612 79736
rect 173020 79868 173084 79932
rect 175228 79868 175292 79932
rect 174860 79792 174924 79796
rect 174860 79736 174874 79792
rect 174874 79736 174924 79792
rect 174860 79732 174924 79736
rect 177252 79792 177316 79796
rect 177252 79736 177256 79792
rect 177256 79736 177312 79792
rect 177312 79736 177316 79792
rect 177252 79732 177316 79736
rect 162716 79460 162780 79524
rect 176700 79460 176764 79524
rect 174676 79384 174740 79388
rect 174676 79328 174726 79384
rect 174726 79328 174740 79384
rect 174676 79324 174740 79328
rect 176516 79324 176580 79388
rect 184796 79188 184860 79252
rect 139900 79052 139964 79116
rect 142660 79052 142724 79116
rect 167868 78976 167932 78980
rect 167868 78920 167882 78976
rect 167882 78920 167932 78976
rect 167868 78916 167932 78920
rect 168236 78976 168300 78980
rect 168236 78920 168286 78976
rect 168286 78920 168300 78976
rect 168236 78916 168300 78920
rect 170812 78976 170876 78980
rect 170812 78920 170862 78976
rect 170862 78920 170876 78976
rect 170812 78916 170876 78920
rect 167132 78780 167196 78844
rect 167868 78780 167932 78844
rect 99236 78644 99300 78708
rect 154068 78644 154132 78708
rect 156092 78644 156156 78708
rect 161244 78644 161308 78708
rect 163452 78644 163516 78708
rect 119292 78508 119356 78572
rect 122236 78568 122300 78572
rect 122236 78512 122286 78568
rect 122286 78512 122300 78568
rect 122236 78508 122300 78512
rect 100340 78372 100404 78436
rect 134932 78508 134996 78572
rect 140452 78508 140516 78572
rect 156644 78568 156708 78572
rect 156644 78512 156658 78568
rect 156658 78512 156708 78568
rect 156644 78508 156708 78512
rect 159588 78508 159652 78572
rect 164924 78508 164988 78572
rect 171732 78508 171796 78572
rect 123892 78372 123956 78436
rect 135668 78372 135732 78436
rect 142108 78372 142172 78436
rect 149284 78372 149348 78436
rect 100524 78236 100588 78300
rect 147996 78236 148060 78300
rect 150940 78236 151004 78300
rect 165844 78236 165908 78300
rect 187004 78372 187068 78436
rect 124076 78100 124140 78164
rect 141188 78160 141252 78164
rect 141188 78104 141238 78160
rect 141238 78104 141252 78160
rect 141188 78100 141252 78104
rect 144500 78100 144564 78164
rect 161980 78100 162044 78164
rect 173020 78160 173084 78164
rect 173020 78104 173070 78160
rect 173070 78104 173084 78160
rect 173020 78100 173084 78104
rect 121132 77964 121196 78028
rect 139348 77964 139412 78028
rect 146708 77964 146772 78028
rect 149284 77964 149348 78028
rect 149652 77964 149716 78028
rect 153700 77964 153764 78028
rect 175044 77964 175108 78028
rect 189212 78100 189276 78164
rect 189028 77964 189092 78028
rect 107148 77692 107212 77756
rect 143580 77828 143644 77892
rect 152780 77828 152844 77892
rect 170812 77828 170876 77892
rect 135852 77692 135916 77756
rect 144132 77692 144196 77756
rect 120948 77556 121012 77620
rect 138244 77556 138308 77620
rect 162900 77556 162964 77620
rect 160692 77148 160756 77212
rect 170812 76876 170876 76940
rect 108436 76740 108500 76804
rect 140268 76800 140332 76804
rect 140268 76744 140282 76800
rect 140282 76744 140332 76800
rect 140268 76740 140332 76744
rect 119844 76604 119908 76668
rect 158116 76664 158180 76668
rect 158116 76608 158130 76664
rect 158130 76608 158180 76664
rect 158116 76604 158180 76608
rect 158300 76604 158364 76668
rect 198780 76604 198844 76668
rect 210372 76740 210436 76804
rect 211108 76604 211172 76668
rect 115428 76468 115492 76532
rect 140084 76332 140148 76396
rect 148548 76196 148612 76260
rect 136220 76060 136284 76124
rect 170628 76060 170692 76124
rect 133092 75924 133156 75988
rect 136404 75984 136468 75988
rect 136404 75928 136418 75984
rect 136418 75928 136468 75984
rect 136404 75924 136468 75928
rect 158852 75984 158916 75988
rect 158852 75928 158866 75984
rect 158866 75928 158916 75984
rect 158852 75924 158916 75928
rect 160508 75984 160572 75988
rect 160508 75928 160522 75984
rect 160522 75928 160572 75984
rect 160508 75924 160572 75928
rect 170076 75984 170140 75988
rect 170076 75928 170090 75984
rect 170090 75928 170140 75984
rect 170076 75924 170140 75928
rect 172284 75924 172348 75988
rect 163452 75788 163516 75852
rect 143948 75652 144012 75716
rect 140636 75380 140700 75444
rect 214052 75380 214116 75444
rect 117084 75244 117148 75308
rect 146708 75244 146772 75308
rect 114140 75108 114204 75172
rect 162348 74428 162412 74492
rect 118372 74292 118436 74356
rect 152596 74292 152660 74356
rect 174676 74292 174740 74356
rect 156092 74156 156156 74220
rect 190500 74156 190564 74220
rect 118188 74020 118252 74084
rect 163636 74020 163700 74084
rect 196204 74020 196268 74084
rect 140452 73884 140516 73948
rect 171732 73884 171796 73948
rect 115612 73748 115676 73812
rect 193628 73748 193692 73812
rect 113036 73612 113100 73676
rect 161796 73612 161860 73676
rect 194732 73612 194796 73676
rect 116716 73068 116780 73132
rect 118556 73128 118620 73132
rect 118556 73072 118570 73128
rect 118570 73072 118620 73128
rect 118556 73068 118620 73072
rect 151124 73068 151188 73132
rect 156644 73128 156708 73132
rect 156644 73072 156658 73128
rect 156658 73072 156708 73128
rect 156644 73068 156708 73072
rect 197308 73068 197372 73132
rect 111012 72932 111076 72996
rect 142660 72796 142724 72860
rect 113588 72524 113652 72588
rect 115796 72388 115860 72452
rect 113956 72252 114020 72316
rect 139348 72252 139412 72316
rect 201540 72796 201604 72860
rect 158484 72660 158548 72724
rect 164556 72524 164620 72588
rect 191972 72388 192036 72452
rect 149652 71708 149716 71772
rect 187188 71708 187252 71772
rect 193444 71572 193508 71636
rect 112668 71436 112732 71500
rect 167684 71436 167748 71500
rect 207612 71436 207676 71500
rect 102916 71300 102980 71364
rect 136588 71300 136652 71364
rect 171548 71300 171612 71364
rect 205588 71300 205652 71364
rect 149284 71164 149348 71228
rect 205772 71164 205836 71228
rect 188108 71028 188172 71092
rect 133092 70892 133156 70956
rect 162900 70892 162964 70956
rect 142108 70408 142172 70412
rect 142108 70352 142122 70408
rect 142122 70352 142172 70408
rect 142108 70348 142172 70352
rect 122604 70212 122668 70276
rect 165844 70212 165908 70276
rect 202092 70212 202156 70276
rect 205036 70212 205100 70276
rect 113772 70076 113836 70140
rect 175044 70076 175108 70140
rect 207060 70076 207124 70140
rect 104572 69940 104636 70004
rect 170628 69940 170692 70004
rect 206140 69940 206204 70004
rect 135300 69804 135364 69868
rect 154252 69804 154316 69868
rect 187740 69804 187804 69868
rect 112852 69668 112916 69732
rect 145052 69668 145116 69732
rect 196572 69668 196636 69732
rect 108804 69532 108868 69596
rect 139900 69532 139964 69596
rect 158300 69532 158364 69596
rect 108620 69396 108684 69460
rect 187924 69396 187988 69460
rect 121316 68852 121380 68916
rect 106964 68716 107028 68780
rect 107332 68580 107396 68644
rect 203012 68580 203076 68644
rect 111564 68444 111628 68508
rect 143580 68444 143644 68508
rect 176516 68444 176580 68508
rect 209820 68444 209884 68508
rect 187372 67492 187436 67556
rect 103284 67356 103348 67420
rect 138244 67356 138308 67420
rect 198964 67356 199028 67420
rect 166580 67220 166644 67284
rect 106044 67084 106108 67148
rect 135852 67084 135916 67148
rect 167868 67084 167932 67148
rect 122972 66948 123036 67012
rect 162716 66948 162780 67012
rect 200620 66948 200684 67012
rect 170996 66812 171060 66876
rect 192156 66676 192220 66740
rect 103100 66132 103164 66196
rect 161060 66132 161124 66196
rect 107516 65996 107580 66060
rect 160692 65996 160756 66060
rect 104756 65860 104820 65924
rect 138060 65860 138124 65924
rect 158116 65860 158180 65924
rect 108252 65724 108316 65788
rect 161980 65724 162044 65788
rect 164924 65588 164988 65652
rect 186084 65452 186148 65516
rect 154436 65316 154500 65380
rect 144132 64772 144196 64836
rect 193260 64772 193324 64836
rect 116900 64636 116964 64700
rect 169156 64636 169220 64700
rect 163452 64500 163516 64564
rect 194548 64500 194612 64564
rect 119660 64364 119724 64428
rect 147812 64364 147876 64428
rect 122052 64228 122116 64292
rect 147996 64228 148060 64292
rect 134932 63820 134996 63884
rect 161244 63412 161308 63476
rect 166764 63276 166828 63340
rect 168052 63140 168116 63204
rect 134932 62052 134996 62116
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 99235 194036 99301 194037
rect 99235 193972 99236 194036
rect 99300 193972 99301 194036
rect 99235 193971 99301 193972
rect 99051 179484 99117 179485
rect 99051 179420 99052 179484
rect 99116 179420 99117 179484
rect 99051 179419 99117 179420
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 99054 80749 99114 179419
rect 99051 80748 99117 80749
rect 99051 80684 99052 80748
rect 99116 80684 99117 80748
rect 99051 80683 99117 80684
rect 99238 78709 99298 193971
rect 100523 180980 100589 180981
rect 100523 180916 100524 180980
rect 100588 180916 100589 180980
rect 100523 180915 100589 180916
rect 100339 148612 100405 148613
rect 100339 148548 100340 148612
rect 100404 148548 100405 148612
rect 100339 148547 100405 148548
rect 99235 78708 99301 78709
rect 99235 78644 99236 78708
rect 99300 78644 99301 78708
rect 99235 78643 99301 78644
rect 100342 78437 100402 148547
rect 100339 78436 100405 78437
rect 100339 78372 100340 78436
rect 100404 78372 100405 78436
rect 100339 78371 100405 78372
rect 100526 78301 100586 180915
rect 100794 174454 101414 209898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 104571 180844 104637 180845
rect 104571 180780 104572 180844
rect 104636 180780 104637 180844
rect 104571 180779 104637 180780
rect 103283 179620 103349 179621
rect 103283 179556 103284 179620
rect 103348 179556 103349 179620
rect 103283 179555 103349 179556
rect 102915 176356 102981 176357
rect 102915 176292 102916 176356
rect 102980 176292 102981 176356
rect 102915 176291 102981 176292
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100523 78300 100589 78301
rect 100523 78236 100524 78300
rect 100588 78236 100589 78300
rect 100523 78235 100589 78236
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 101898
rect 102918 71365 102978 176291
rect 103099 176220 103165 176221
rect 103099 176156 103100 176220
rect 103164 176156 103165 176220
rect 103099 176155 103165 176156
rect 102915 71364 102981 71365
rect 102915 71300 102916 71364
rect 102980 71300 102981 71364
rect 102915 71299 102981 71300
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 103102 66197 103162 176155
rect 103286 67421 103346 179555
rect 104574 70005 104634 180779
rect 104755 180164 104821 180165
rect 104755 180100 104756 180164
rect 104820 180100 104821 180164
rect 104755 180099 104821 180100
rect 104571 70004 104637 70005
rect 104571 69940 104572 70004
rect 104636 69940 104637 70004
rect 104571 69939 104637 69940
rect 103283 67420 103349 67421
rect 103283 67356 103284 67420
rect 103348 67356 103349 67420
rect 103283 67355 103349 67356
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 103099 66196 103165 66197
rect 103099 66132 103100 66196
rect 103164 66132 103165 66196
rect 103099 66131 103165 66132
rect 104758 65925 104818 180099
rect 105294 178954 105914 214398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 111747 265572 111813 265573
rect 111747 265508 111748 265572
rect 111812 265508 111813 265572
rect 111747 265507 111813 265508
rect 111750 262853 111810 265507
rect 111747 262852 111813 262853
rect 111747 262788 111748 262852
rect 111812 262788 111813 262852
rect 111747 262787 111813 262788
rect 112851 262852 112917 262853
rect 112851 262788 112852 262852
rect 112916 262788 112917 262852
rect 112851 262787 112917 262788
rect 111563 259724 111629 259725
rect 111563 259660 111564 259724
rect 111628 259660 111629 259724
rect 111563 259659 111629 259660
rect 111379 259588 111445 259589
rect 111379 259524 111380 259588
rect 111444 259524 111445 259588
rect 111379 259523 111445 259524
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 107515 199476 107581 199477
rect 107515 199412 107516 199476
rect 107580 199412 107581 199476
rect 107515 199411 107581 199412
rect 107518 198797 107578 199411
rect 107515 198796 107581 198797
rect 107515 198732 107516 198796
rect 107580 198732 107581 198796
rect 107515 198731 107581 198732
rect 107147 182884 107213 182885
rect 107147 182820 107148 182884
rect 107212 182820 107213 182884
rect 107147 182819 107213 182820
rect 106043 179756 106109 179757
rect 106043 179692 106044 179756
rect 106108 179692 106109 179756
rect 106043 179691 106109 179692
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 100794 30454 101414 65898
rect 104755 65924 104821 65925
rect 104755 65860 104756 65924
rect 104820 65860 104821 65924
rect 104755 65859 104821 65860
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 70398
rect 106046 67149 106106 179691
rect 106963 148340 107029 148341
rect 106963 148276 106964 148340
rect 107028 148276 107029 148340
rect 106963 148275 107029 148276
rect 106966 68781 107026 148275
rect 107150 77757 107210 182819
rect 107331 180028 107397 180029
rect 107331 179964 107332 180028
rect 107396 179964 107397 180028
rect 107331 179963 107397 179964
rect 107147 77756 107213 77757
rect 107147 77692 107148 77756
rect 107212 77692 107213 77756
rect 107147 77691 107213 77692
rect 106963 68780 107029 68781
rect 106963 68716 106964 68780
rect 107028 68716 107029 68780
rect 106963 68715 107029 68716
rect 107334 68645 107394 179963
rect 107331 68644 107397 68645
rect 107331 68580 107332 68644
rect 107396 68580 107397 68644
rect 107331 68579 107397 68580
rect 106043 67148 106109 67149
rect 106043 67084 106044 67148
rect 106108 67084 106109 67148
rect 106043 67083 106109 67084
rect 107518 66061 107578 198731
rect 108803 194172 108869 194173
rect 108803 194108 108804 194172
rect 108868 194108 108869 194172
rect 108803 194107 108869 194108
rect 108435 187100 108501 187101
rect 108435 187036 108436 187100
rect 108500 187036 108501 187100
rect 108435 187035 108501 187036
rect 108251 138820 108317 138821
rect 108251 138756 108252 138820
rect 108316 138756 108317 138820
rect 108251 138755 108317 138756
rect 107515 66060 107581 66061
rect 107515 65996 107516 66060
rect 107580 65996 107581 66060
rect 107515 65995 107581 65996
rect 108254 65789 108314 138755
rect 108438 76805 108498 187035
rect 108619 182204 108685 182205
rect 108619 182140 108620 182204
rect 108684 182140 108685 182204
rect 108619 182139 108685 182140
rect 108435 76804 108501 76805
rect 108435 76740 108436 76804
rect 108500 76740 108501 76804
rect 108435 76739 108501 76740
rect 108622 69461 108682 182139
rect 108806 69597 108866 194107
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 111011 148476 111077 148477
rect 111011 148412 111012 148476
rect 111076 148412 111077 148476
rect 111011 148411 111077 148412
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 108803 69596 108869 69597
rect 108803 69532 108804 69596
rect 108868 69532 108869 69596
rect 108803 69531 108869 69532
rect 108619 69460 108685 69461
rect 108619 69396 108620 69460
rect 108684 69396 108685 69460
rect 108619 69395 108685 69396
rect 108251 65788 108317 65789
rect 108251 65724 108252 65788
rect 108316 65724 108317 65788
rect 108251 65723 108317 65724
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 74898
rect 111014 72997 111074 148411
rect 111382 145893 111442 259523
rect 111566 146029 111626 259659
rect 112483 186964 112549 186965
rect 112483 186900 112484 186964
rect 112548 186900 112549 186964
rect 112483 186899 112549 186900
rect 111563 146028 111629 146029
rect 111563 145964 111564 146028
rect 111628 145964 111629 146028
rect 111563 145963 111629 145964
rect 111379 145892 111445 145893
rect 111379 145828 111380 145892
rect 111444 145828 111445 145892
rect 111379 145827 111445 145828
rect 111563 144396 111629 144397
rect 111563 144332 111564 144396
rect 111628 144332 111629 144396
rect 111563 144331 111629 144332
rect 111195 137868 111261 137869
rect 111195 137804 111196 137868
rect 111260 137804 111261 137868
rect 111195 137803 111261 137804
rect 111198 81701 111258 137803
rect 111195 81700 111261 81701
rect 111195 81636 111196 81700
rect 111260 81636 111261 81700
rect 111195 81635 111261 81636
rect 111011 72996 111077 72997
rect 111011 72932 111012 72996
rect 111076 72932 111077 72996
rect 111011 72931 111077 72932
rect 111566 68509 111626 144331
rect 112486 80885 112546 186899
rect 112667 185604 112733 185605
rect 112667 185540 112668 185604
rect 112732 185540 112733 185604
rect 112667 185539 112733 185540
rect 112483 80884 112549 80885
rect 112483 80820 112484 80884
rect 112548 80820 112549 80884
rect 112483 80819 112549 80820
rect 112670 71501 112730 185539
rect 112854 145757 112914 262787
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118555 263940 118621 263941
rect 118555 263876 118556 263940
rect 118620 263876 118621 263940
rect 118555 263875 118621 263876
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 116899 263804 116965 263805
rect 116899 263740 116900 263804
rect 116964 263740 116965 263804
rect 116899 263739 116965 263740
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114139 191044 114205 191045
rect 114139 190980 114140 191044
rect 114204 190980 114205 191044
rect 114139 190979 114205 190980
rect 113035 190500 113101 190501
rect 113035 190436 113036 190500
rect 113100 190436 113101 190500
rect 113035 190435 113101 190436
rect 112851 145756 112917 145757
rect 112851 145692 112852 145756
rect 112916 145692 112917 145756
rect 112851 145691 112917 145692
rect 112851 141948 112917 141949
rect 112851 141884 112852 141948
rect 112916 141884 112917 141948
rect 112851 141883 112917 141884
rect 112667 71500 112733 71501
rect 112667 71436 112668 71500
rect 112732 71436 112733 71500
rect 112667 71435 112733 71436
rect 112854 69733 112914 141883
rect 113038 73677 113098 190435
rect 113955 187236 114021 187237
rect 113955 187172 113956 187236
rect 114020 187172 114021 187236
rect 113955 187171 114021 187172
rect 113771 144124 113837 144125
rect 113771 144060 113772 144124
rect 113836 144060 113837 144124
rect 113771 144059 113837 144060
rect 113587 140452 113653 140453
rect 113587 140388 113588 140452
rect 113652 140388 113653 140452
rect 113587 140387 113653 140388
rect 113035 73676 113101 73677
rect 113035 73612 113036 73676
rect 113100 73612 113101 73676
rect 113035 73611 113101 73612
rect 113590 72589 113650 140387
rect 113587 72588 113653 72589
rect 113587 72524 113588 72588
rect 113652 72524 113653 72588
rect 113587 72523 113653 72524
rect 113774 70141 113834 144059
rect 113958 72317 114018 187171
rect 114142 75173 114202 190979
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 116531 144260 116597 144261
rect 116531 144196 116532 144260
rect 116596 144196 116597 144260
rect 116531 144195 116597 144196
rect 115611 140588 115677 140589
rect 115611 140524 115612 140588
rect 115676 140524 115677 140588
rect 115611 140523 115677 140524
rect 115427 139908 115493 139909
rect 115427 139844 115428 139908
rect 115492 139844 115493 139908
rect 115427 139843 115493 139844
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114139 75172 114205 75173
rect 114139 75108 114140 75172
rect 114204 75108 114205 75172
rect 114139 75107 114205 75108
rect 113955 72316 114021 72317
rect 113955 72252 113956 72316
rect 114020 72252 114021 72316
rect 113955 72251 114021 72252
rect 113771 70140 113837 70141
rect 113771 70076 113772 70140
rect 113836 70076 113837 70140
rect 113771 70075 113837 70076
rect 112851 69732 112917 69733
rect 112851 69668 112852 69732
rect 112916 69668 112917 69732
rect 112851 69667 112917 69668
rect 111563 68508 111629 68509
rect 111563 68444 111564 68508
rect 111628 68444 111629 68508
rect 111563 68443 111629 68444
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 79398
rect 115430 76533 115490 139843
rect 115427 76532 115493 76533
rect 115427 76468 115428 76532
rect 115492 76468 115493 76532
rect 115427 76467 115493 76468
rect 115614 73813 115674 140523
rect 115795 138140 115861 138141
rect 115795 138076 115796 138140
rect 115860 138076 115861 138140
rect 115795 138075 115861 138076
rect 115611 73812 115677 73813
rect 115611 73748 115612 73812
rect 115676 73748 115677 73812
rect 115611 73747 115677 73748
rect 115798 72453 115858 138075
rect 116534 80613 116594 144195
rect 116902 143037 116962 263739
rect 117083 196620 117149 196621
rect 117083 196556 117084 196620
rect 117148 196556 117149 196620
rect 117083 196555 117149 196556
rect 116899 143036 116965 143037
rect 116899 142972 116900 143036
rect 116964 142972 116965 143036
rect 116899 142971 116965 142972
rect 116715 141404 116781 141405
rect 116715 141340 116716 141404
rect 116780 141340 116781 141404
rect 116715 141339 116781 141340
rect 116531 80612 116597 80613
rect 116531 80548 116532 80612
rect 116596 80548 116597 80612
rect 116531 80547 116597 80548
rect 116718 73133 116778 141339
rect 116899 139500 116965 139501
rect 116899 139436 116900 139500
rect 116964 139436 116965 139500
rect 116899 139435 116965 139436
rect 116715 73132 116781 73133
rect 116715 73068 116716 73132
rect 116780 73068 116781 73132
rect 116715 73067 116781 73068
rect 115795 72452 115861 72453
rect 115795 72388 115796 72452
rect 115860 72388 115861 72452
rect 115795 72387 115861 72388
rect 116902 64701 116962 139435
rect 117086 75309 117146 196555
rect 118371 189684 118437 189685
rect 118371 189620 118372 189684
rect 118436 189620 118437 189684
rect 118371 189619 118437 189620
rect 118187 141540 118253 141541
rect 118187 141476 118188 141540
rect 118252 141476 118253 141540
rect 118187 141475 118253 141476
rect 117083 75308 117149 75309
rect 117083 75244 117084 75308
rect 117148 75244 117149 75308
rect 117083 75243 117149 75244
rect 118190 74085 118250 141475
rect 118374 74357 118434 189619
rect 118558 142901 118618 263875
rect 118794 262000 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 121499 262308 121565 262309
rect 121499 262244 121500 262308
rect 121564 262244 121565 262308
rect 121499 262243 121565 262244
rect 121315 260132 121381 260133
rect 121315 260068 121316 260132
rect 121380 260068 121381 260132
rect 121315 260067 121381 260068
rect 118794 192454 119414 198000
rect 121318 194581 121378 260067
rect 121502 218109 121562 262243
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 196019 269788 196085 269789
rect 196019 269724 196020 269788
rect 196084 269724 196085 269788
rect 196019 269723 196085 269724
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 194547 268428 194613 268429
rect 194547 268364 194548 268428
rect 194612 268364 194613 268428
rect 194547 268363 194613 268364
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 262000 191414 263898
rect 191787 262988 191853 262989
rect 191787 262924 191788 262988
rect 191852 262924 191853 262988
rect 191787 262923 191853 262924
rect 122603 259996 122669 259997
rect 122603 259932 122604 259996
rect 122668 259932 122669 259996
rect 122603 259931 122669 259932
rect 187187 259996 187253 259997
rect 187187 259932 187188 259996
rect 187252 259932 187253 259996
rect 187187 259931 187253 259932
rect 122051 237420 122117 237421
rect 122051 237356 122052 237420
rect 122116 237356 122117 237420
rect 122051 237355 122117 237356
rect 121499 218108 121565 218109
rect 121499 218044 121500 218108
rect 121564 218044 121565 218108
rect 121499 218043 121565 218044
rect 122054 200429 122114 237355
rect 122235 216748 122301 216749
rect 122235 216684 122236 216748
rect 122300 216684 122301 216748
rect 122235 216683 122301 216684
rect 122238 200837 122298 216683
rect 122419 212668 122485 212669
rect 122419 212604 122420 212668
rect 122484 212604 122485 212668
rect 122419 212603 122485 212604
rect 122235 200836 122301 200837
rect 122235 200772 122236 200836
rect 122300 200772 122301 200836
rect 122235 200771 122301 200772
rect 122051 200428 122117 200429
rect 122051 200364 122052 200428
rect 122116 200364 122117 200428
rect 122051 200363 122117 200364
rect 122422 199477 122482 212603
rect 122419 199476 122485 199477
rect 122419 199412 122420 199476
rect 122484 199412 122485 199476
rect 122419 199411 122485 199412
rect 122235 196756 122301 196757
rect 122235 196692 122236 196756
rect 122300 196692 122301 196756
rect 122235 196691 122301 196692
rect 121315 194580 121381 194581
rect 121315 194516 121316 194580
rect 121380 194516 121381 194580
rect 121315 194515 121381 194516
rect 119659 193900 119725 193901
rect 119659 193836 119660 193900
rect 119724 193836 119725 193900
rect 119659 193835 119725 193836
rect 119662 192949 119722 193835
rect 119659 192948 119725 192949
rect 119659 192884 119660 192948
rect 119724 192884 119725 192948
rect 119659 192883 119725 192884
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 119662 190470 119722 192883
rect 119662 190410 119906 190470
rect 119659 189820 119725 189821
rect 119659 189756 119660 189820
rect 119724 189756 119725 189820
rect 119659 189755 119725 189756
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118555 142900 118621 142901
rect 118555 142836 118556 142900
rect 118620 142836 118621 142900
rect 118555 142835 118621 142836
rect 118794 142000 119414 155898
rect 118555 141676 118621 141677
rect 118555 141612 118556 141676
rect 118620 141612 118621 141676
rect 118555 141611 118621 141612
rect 118371 74356 118437 74357
rect 118371 74292 118372 74356
rect 118436 74292 118437 74356
rect 118371 74291 118437 74292
rect 118187 74084 118253 74085
rect 118187 74020 118188 74084
rect 118252 74020 118253 74084
rect 118187 74019 118253 74020
rect 118558 73133 118618 141611
rect 119662 89730 119722 189755
rect 119294 89670 119722 89730
rect 119294 78573 119354 89670
rect 119659 81564 119725 81565
rect 119659 81500 119660 81564
rect 119724 81500 119725 81564
rect 119659 81499 119725 81500
rect 119291 78572 119357 78573
rect 119291 78508 119292 78572
rect 119356 78508 119357 78572
rect 119291 78507 119357 78508
rect 118555 73132 118621 73133
rect 118555 73068 118556 73132
rect 118620 73068 118621 73132
rect 118555 73067 118621 73068
rect 116899 64700 116965 64701
rect 116899 64636 116900 64700
rect 116964 64636 116965 64700
rect 116899 64635 116965 64636
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 119662 64429 119722 81499
rect 119846 76669 119906 190410
rect 122238 176629 122298 196691
rect 122606 195941 122666 259931
rect 187003 259316 187069 259317
rect 187003 259252 187004 259316
rect 187068 259252 187069 259316
rect 187003 259251 187069 259252
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 186819 233340 186885 233341
rect 186819 233276 186820 233340
rect 186884 233276 186885 233340
rect 186819 233275 186885 233276
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 181483 201788 181549 201789
rect 181483 201724 181484 201788
rect 181548 201724 181549 201788
rect 181483 201723 181549 201724
rect 138611 201516 138677 201517
rect 138611 201452 138612 201516
rect 138676 201452 138677 201516
rect 138611 201451 138677 201452
rect 160323 201516 160389 201517
rect 160323 201452 160324 201516
rect 160388 201452 160389 201516
rect 160323 201451 160389 201452
rect 137875 200700 137941 200701
rect 137875 200636 137876 200700
rect 137940 200636 137941 200700
rect 137875 200635 137941 200636
rect 133643 199884 133709 199885
rect 133643 199820 133644 199884
rect 133708 199820 133709 199884
rect 133643 199819 133709 199820
rect 133827 199884 133893 199885
rect 133827 199820 133828 199884
rect 133892 199820 133893 199884
rect 133827 199819 133893 199820
rect 134195 199884 134261 199885
rect 134195 199820 134196 199884
rect 134260 199820 134261 199884
rect 134195 199819 134261 199820
rect 135115 199884 135181 199885
rect 135115 199820 135116 199884
rect 135180 199820 135181 199884
rect 135115 199819 135181 199820
rect 136219 199884 136285 199885
rect 136219 199820 136220 199884
rect 136284 199820 136285 199884
rect 136219 199819 136285 199820
rect 123294 196954 123914 198000
rect 133646 197165 133706 199819
rect 132539 197164 132605 197165
rect 132539 197100 132540 197164
rect 132604 197100 132605 197164
rect 132539 197099 132605 197100
rect 133643 197164 133709 197165
rect 133643 197100 133644 197164
rect 133708 197100 133709 197164
rect 133643 197099 133709 197100
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122603 195940 122669 195941
rect 122603 195876 122604 195940
rect 122668 195876 122669 195940
rect 122603 195875 122669 195876
rect 122603 191180 122669 191181
rect 122603 191116 122604 191180
rect 122668 191116 122669 191180
rect 122603 191115 122669 191116
rect 122419 188596 122485 188597
rect 122419 188532 122420 188596
rect 122484 188532 122485 188596
rect 122419 188531 122485 188532
rect 122235 176628 122301 176629
rect 122235 176564 122236 176628
rect 122300 176564 122301 176628
rect 122235 176563 122301 176564
rect 121131 176492 121197 176493
rect 121131 176428 121132 176492
rect 121196 176428 121197 176492
rect 121131 176427 121197 176428
rect 120947 140724 121013 140725
rect 120947 140660 120948 140724
rect 121012 140660 121013 140724
rect 120947 140659 121013 140660
rect 120579 140180 120645 140181
rect 120579 140116 120580 140180
rect 120644 140116 120645 140180
rect 120579 140115 120645 140116
rect 120582 92581 120642 140115
rect 120579 92580 120645 92581
rect 120579 92516 120580 92580
rect 120644 92516 120645 92580
rect 120579 92515 120645 92516
rect 120950 77621 121010 140659
rect 121134 78029 121194 176427
rect 121315 175948 121381 175949
rect 121315 175884 121316 175948
rect 121380 175884 121381 175948
rect 121315 175883 121381 175884
rect 121131 78028 121197 78029
rect 121131 77964 121132 78028
rect 121196 77964 121197 78028
rect 121131 77963 121197 77964
rect 120947 77620 121013 77621
rect 120947 77556 120948 77620
rect 121012 77556 121013 77620
rect 120947 77555 121013 77556
rect 119843 76668 119909 76669
rect 119843 76604 119844 76668
rect 119908 76604 119909 76668
rect 119843 76603 119909 76604
rect 121318 68917 121378 175883
rect 121867 140044 121933 140045
rect 121867 139980 121868 140044
rect 121932 139980 121933 140044
rect 121867 139979 121933 139980
rect 121870 122850 121930 139979
rect 122051 139364 122117 139365
rect 122051 139300 122052 139364
rect 122116 139300 122117 139364
rect 122051 139299 122117 139300
rect 122054 132701 122114 139299
rect 122051 132700 122117 132701
rect 122051 132636 122052 132700
rect 122116 132636 122117 132700
rect 122051 132635 122117 132636
rect 122051 132428 122117 132429
rect 122051 132364 122052 132428
rect 122116 132364 122117 132428
rect 122051 132363 122117 132364
rect 122054 123045 122114 132363
rect 122051 123044 122117 123045
rect 122051 122980 122052 123044
rect 122116 122980 122117 123044
rect 122051 122979 122117 122980
rect 121870 122790 122114 122850
rect 121315 68916 121381 68917
rect 121315 68852 121316 68916
rect 121380 68852 121381 68916
rect 121315 68851 121381 68852
rect 119659 64428 119725 64429
rect 119659 64364 119660 64428
rect 119724 64364 119725 64428
rect 119659 64363 119725 64364
rect 122054 64293 122114 122790
rect 122238 78573 122298 176563
rect 122422 79389 122482 188531
rect 122419 79388 122485 79389
rect 122419 79324 122420 79388
rect 122484 79324 122485 79388
rect 122419 79323 122485 79324
rect 122235 78572 122301 78573
rect 122235 78508 122236 78572
rect 122300 78508 122301 78572
rect 122235 78507 122301 78508
rect 122606 70277 122666 191115
rect 122971 187372 123037 187373
rect 122971 187308 122972 187372
rect 123036 187308 123037 187372
rect 122971 187307 123037 187308
rect 122974 138005 123034 187307
rect 123294 160954 123914 196398
rect 124075 195668 124141 195669
rect 124075 195604 124076 195668
rect 124140 195604 124141 195668
rect 124075 195603 124141 195604
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 123891 139364 123957 139365
rect 123891 139300 123892 139364
rect 123956 139300 123957 139364
rect 123891 139299 123957 139300
rect 122971 138004 123037 138005
rect 122971 137940 122972 138004
rect 123036 137940 123037 138004
rect 122971 137939 123037 137940
rect 122787 132700 122853 132701
rect 122787 132636 122788 132700
rect 122852 132636 122853 132700
rect 122787 132635 122853 132636
rect 122790 132429 122850 132635
rect 122787 132428 122853 132429
rect 122787 132364 122788 132428
rect 122852 132364 122853 132428
rect 122787 132363 122853 132364
rect 122787 123044 122853 123045
rect 122787 122980 122788 123044
rect 122852 122980 122853 123044
rect 122787 122979 122853 122980
rect 122790 122773 122850 122979
rect 122787 122772 122853 122773
rect 122787 122708 122788 122772
rect 122852 122708 122853 122772
rect 122787 122707 122853 122708
rect 122787 113252 122853 113253
rect 122787 113188 122788 113252
rect 122852 113188 122853 113252
rect 122787 113187 122853 113188
rect 122790 113117 122850 113187
rect 122787 113116 122853 113117
rect 122787 113052 122788 113116
rect 122852 113052 122853 113116
rect 122787 113051 122853 113052
rect 122787 103596 122853 103597
rect 122787 103532 122788 103596
rect 122852 103532 122853 103596
rect 122787 103531 122853 103532
rect 122790 103461 122850 103531
rect 122787 103460 122853 103461
rect 122787 103396 122788 103460
rect 122852 103396 122853 103460
rect 122787 103395 122853 103396
rect 122787 93940 122853 93941
rect 122787 93876 122788 93940
rect 122852 93876 122853 93940
rect 122787 93875 122853 93876
rect 122790 93805 122850 93875
rect 122787 93804 122853 93805
rect 122787 93740 122788 93804
rect 122852 93740 122853 93804
rect 122787 93739 122853 93740
rect 122971 83468 123037 83469
rect 122971 83404 122972 83468
rect 123036 83404 123037 83468
rect 122971 83403 123037 83404
rect 122603 70276 122669 70277
rect 122603 70212 122604 70276
rect 122668 70212 122669 70276
rect 122603 70211 122669 70212
rect 122974 67013 123034 83403
rect 123894 78437 123954 139299
rect 123891 78436 123957 78437
rect 123891 78372 123892 78436
rect 123956 78372 123957 78436
rect 123891 78371 123957 78372
rect 124078 78165 124138 195603
rect 132542 188461 132602 197099
rect 133830 196485 133890 199819
rect 133827 196484 133893 196485
rect 133827 196420 133828 196484
rect 133892 196420 133893 196484
rect 133827 196419 133893 196420
rect 134198 193357 134258 199819
rect 134379 197844 134445 197845
rect 134379 197780 134380 197844
rect 134444 197780 134445 197844
rect 134379 197779 134445 197780
rect 134195 193356 134261 193357
rect 134195 193292 134196 193356
rect 134260 193292 134261 193356
rect 134195 193291 134261 193292
rect 132539 188460 132605 188461
rect 132539 188396 132540 188460
rect 132604 188396 132605 188460
rect 132539 188395 132605 188396
rect 124811 176084 124877 176085
rect 124811 176020 124812 176084
rect 124876 176020 124877 176084
rect 124811 176019 124877 176020
rect 124814 137869 124874 176019
rect 134382 140317 134442 197779
rect 135118 196349 135178 199819
rect 135851 199612 135917 199613
rect 135851 199548 135852 199612
rect 135916 199548 135917 199612
rect 135851 199547 135917 199548
rect 135115 196348 135181 196349
rect 135115 196284 135116 196348
rect 135180 196284 135181 196348
rect 135115 196283 135181 196284
rect 135854 175949 135914 199547
rect 136035 195940 136101 195941
rect 136035 195876 136036 195940
rect 136100 195876 136101 195940
rect 136035 195875 136101 195876
rect 136038 177853 136098 195875
rect 136222 179485 136282 199819
rect 136403 199748 136469 199749
rect 136403 199684 136404 199748
rect 136468 199684 136469 199748
rect 136403 199683 136469 199684
rect 136406 195941 136466 199683
rect 137878 196485 137938 200635
rect 138427 199884 138493 199885
rect 138427 199820 138428 199884
rect 138492 199820 138493 199884
rect 138427 199819 138493 199820
rect 138243 199748 138309 199749
rect 138243 199684 138244 199748
rect 138308 199684 138309 199748
rect 138243 199683 138309 199684
rect 138246 196757 138306 199683
rect 138243 196756 138309 196757
rect 138243 196692 138244 196756
rect 138308 196692 138309 196756
rect 138243 196691 138309 196692
rect 137875 196484 137941 196485
rect 137875 196420 137876 196484
rect 137940 196420 137941 196484
rect 137875 196419 137941 196420
rect 137323 196212 137389 196213
rect 137323 196148 137324 196212
rect 137388 196148 137389 196212
rect 137323 196147 137389 196148
rect 137875 196212 137941 196213
rect 137875 196148 137876 196212
rect 137940 196148 137941 196212
rect 137875 196147 137941 196148
rect 136403 195940 136469 195941
rect 136403 195876 136404 195940
rect 136468 195876 136469 195940
rect 136403 195875 136469 195876
rect 137139 195940 137205 195941
rect 137139 195876 137140 195940
rect 137204 195876 137205 195940
rect 137139 195875 137205 195876
rect 136219 179484 136285 179485
rect 136219 179420 136220 179484
rect 136284 179420 136285 179484
rect 136219 179419 136285 179420
rect 136035 177852 136101 177853
rect 136035 177788 136036 177852
rect 136100 177788 136101 177852
rect 136035 177787 136101 177788
rect 137142 176357 137202 195875
rect 137326 190365 137386 196147
rect 137323 190364 137389 190365
rect 137323 190300 137324 190364
rect 137388 190300 137389 190364
rect 137323 190299 137389 190300
rect 137878 180709 137938 196147
rect 138430 195941 138490 199819
rect 138614 199749 138674 201451
rect 154251 200972 154317 200973
rect 154251 200908 154252 200972
rect 154316 200908 154317 200972
rect 154251 200907 154317 200908
rect 146523 200836 146589 200837
rect 146523 200772 146524 200836
rect 146588 200772 146589 200836
rect 146523 200771 146589 200772
rect 140451 200292 140517 200293
rect 140451 200228 140452 200292
rect 140516 200228 140517 200292
rect 140451 200227 140517 200228
rect 138795 199884 138861 199885
rect 138795 199820 138796 199884
rect 138860 199820 138861 199884
rect 138795 199819 138861 199820
rect 139347 199884 139413 199885
rect 139347 199820 139348 199884
rect 139412 199820 139413 199884
rect 139347 199819 139413 199820
rect 140083 199884 140149 199885
rect 140083 199820 140084 199884
rect 140148 199820 140149 199884
rect 140083 199819 140149 199820
rect 140267 199884 140333 199885
rect 140267 199820 140268 199884
rect 140332 199820 140333 199884
rect 140267 199819 140333 199820
rect 138611 199748 138677 199749
rect 138611 199684 138612 199748
rect 138676 199684 138677 199748
rect 138611 199683 138677 199684
rect 138798 198661 138858 199819
rect 138795 198660 138861 198661
rect 138795 198596 138796 198660
rect 138860 198596 138861 198660
rect 138795 198595 138861 198596
rect 138979 198252 139045 198253
rect 138979 198188 138980 198252
rect 139044 198188 139045 198252
rect 138979 198187 139045 198188
rect 138795 196484 138861 196485
rect 138795 196420 138796 196484
rect 138860 196420 138861 196484
rect 138795 196419 138861 196420
rect 138427 195940 138493 195941
rect 138427 195876 138428 195940
rect 138492 195876 138493 195940
rect 138427 195875 138493 195876
rect 138611 195940 138677 195941
rect 138611 195876 138612 195940
rect 138676 195876 138677 195940
rect 138611 195875 138677 195876
rect 137875 180708 137941 180709
rect 137875 180644 137876 180708
rect 137940 180644 137941 180708
rect 137875 180643 137941 180644
rect 137878 179485 137938 180643
rect 138614 180165 138674 195875
rect 138798 180845 138858 196419
rect 138982 183565 139042 198187
rect 139350 196077 139410 199819
rect 139715 199748 139781 199749
rect 139715 199684 139716 199748
rect 139780 199684 139781 199748
rect 139715 199683 139781 199684
rect 139718 199205 139778 199683
rect 140086 199205 140146 199819
rect 139715 199204 139781 199205
rect 139715 199140 139716 199204
rect 139780 199140 139781 199204
rect 139715 199139 139781 199140
rect 140083 199204 140149 199205
rect 140083 199140 140084 199204
rect 140148 199140 140149 199204
rect 140083 199139 140149 199140
rect 140270 198525 140330 199819
rect 140454 199205 140514 200227
rect 146526 199885 146586 200771
rect 152595 200156 152661 200157
rect 152595 200092 152596 200156
rect 152660 200092 152661 200156
rect 152595 200091 152661 200092
rect 141003 199884 141069 199885
rect 141003 199820 141004 199884
rect 141068 199820 141069 199884
rect 141003 199819 141069 199820
rect 142475 199884 142541 199885
rect 142475 199820 142476 199884
rect 142540 199820 142541 199884
rect 142475 199819 142541 199820
rect 144683 199884 144749 199885
rect 144683 199820 144684 199884
rect 144748 199820 144749 199884
rect 144683 199819 144749 199820
rect 145235 199884 145301 199885
rect 145235 199820 145236 199884
rect 145300 199820 145301 199884
rect 145235 199819 145301 199820
rect 146523 199884 146589 199885
rect 146523 199820 146524 199884
rect 146588 199820 146589 199884
rect 146523 199819 146589 199820
rect 147443 199884 147509 199885
rect 147443 199820 147444 199884
rect 147508 199820 147509 199884
rect 147443 199819 147509 199820
rect 147995 199884 148061 199885
rect 147995 199820 147996 199884
rect 148060 199820 148061 199884
rect 147995 199819 148061 199820
rect 149467 199884 149533 199885
rect 149467 199820 149468 199884
rect 149532 199820 149533 199884
rect 149467 199819 149533 199820
rect 150019 199884 150085 199885
rect 150019 199820 150020 199884
rect 150084 199820 150085 199884
rect 150019 199819 150085 199820
rect 150571 199884 150637 199885
rect 150571 199820 150572 199884
rect 150636 199820 150637 199884
rect 150571 199819 150637 199820
rect 151123 199884 151189 199885
rect 151123 199820 151124 199884
rect 151188 199820 151189 199884
rect 151123 199819 151189 199820
rect 140451 199204 140517 199205
rect 140451 199140 140452 199204
rect 140516 199140 140517 199204
rect 140451 199139 140517 199140
rect 140267 198524 140333 198525
rect 140267 198460 140268 198524
rect 140332 198460 140333 198524
rect 140267 198459 140333 198460
rect 141006 197845 141066 199819
rect 141371 199748 141437 199749
rect 141371 199684 141372 199748
rect 141436 199684 141437 199748
rect 141371 199683 141437 199684
rect 141374 198253 141434 199683
rect 142291 198524 142357 198525
rect 142291 198460 142292 198524
rect 142356 198460 142357 198524
rect 142291 198459 142357 198460
rect 141371 198252 141437 198253
rect 141371 198188 141372 198252
rect 141436 198188 141437 198252
rect 141371 198187 141437 198188
rect 141003 197844 141069 197845
rect 141003 197780 141004 197844
rect 141068 197780 141069 197844
rect 141003 197779 141069 197780
rect 141003 197164 141069 197165
rect 141003 197100 141004 197164
rect 141068 197100 141069 197164
rect 141003 197099 141069 197100
rect 139899 196756 139965 196757
rect 139899 196692 139900 196756
rect 139964 196692 139965 196756
rect 139899 196691 139965 196692
rect 139347 196076 139413 196077
rect 139347 196012 139348 196076
rect 139412 196012 139413 196076
rect 139347 196011 139413 196012
rect 138979 183564 139045 183565
rect 138979 183500 138980 183564
rect 139044 183500 139045 183564
rect 138979 183499 139045 183500
rect 139902 182885 139962 196691
rect 139899 182884 139965 182885
rect 139899 182820 139900 182884
rect 139964 182820 139965 182884
rect 139899 182819 139965 182820
rect 138795 180844 138861 180845
rect 138795 180780 138796 180844
rect 138860 180780 138861 180844
rect 138795 180779 138861 180780
rect 138798 180437 138858 180779
rect 138795 180436 138861 180437
rect 138795 180372 138796 180436
rect 138860 180372 138861 180436
rect 138795 180371 138861 180372
rect 138611 180164 138677 180165
rect 138611 180100 138612 180164
rect 138676 180100 138677 180164
rect 138611 180099 138677 180100
rect 137875 179484 137941 179485
rect 137875 179420 137876 179484
rect 137940 179420 137941 179484
rect 137875 179419 137941 179420
rect 141006 177989 141066 197099
rect 141294 178954 141914 198000
rect 142294 194173 142354 198459
rect 142478 197437 142538 199819
rect 143027 199748 143093 199749
rect 143027 199684 143028 199748
rect 143092 199684 143093 199748
rect 143027 199683 143093 199684
rect 143947 199748 144013 199749
rect 143947 199684 143948 199748
rect 144012 199684 144013 199748
rect 143947 199683 144013 199684
rect 142475 197436 142541 197437
rect 142475 197372 142476 197436
rect 142540 197372 142541 197436
rect 142475 197371 142541 197372
rect 143030 195125 143090 199683
rect 143211 199612 143277 199613
rect 143211 199548 143212 199612
rect 143276 199548 143277 199612
rect 143211 199547 143277 199548
rect 143579 199612 143645 199613
rect 143579 199548 143580 199612
rect 143644 199548 143645 199612
rect 143579 199547 143645 199548
rect 143214 196757 143274 199547
rect 143395 199068 143461 199069
rect 143395 199004 143396 199068
rect 143460 199004 143461 199068
rect 143395 199003 143461 199004
rect 143211 196756 143277 196757
rect 143211 196692 143212 196756
rect 143276 196692 143277 196756
rect 143211 196691 143277 196692
rect 143027 195124 143093 195125
rect 143027 195060 143028 195124
rect 143092 195060 143093 195124
rect 143027 195059 143093 195060
rect 142291 194172 142357 194173
rect 142291 194108 142292 194172
rect 142356 194108 142357 194172
rect 142291 194107 142357 194108
rect 143398 188733 143458 199003
rect 143395 188732 143461 188733
rect 143395 188668 143396 188732
rect 143460 188668 143461 188732
rect 143395 188667 143461 188668
rect 143582 188325 143642 199547
rect 143950 195941 144010 199683
rect 144499 198524 144565 198525
rect 144499 198460 144500 198524
rect 144564 198460 144565 198524
rect 144499 198459 144565 198460
rect 144131 197164 144197 197165
rect 144131 197100 144132 197164
rect 144196 197100 144197 197164
rect 144131 197099 144197 197100
rect 143947 195940 144013 195941
rect 143947 195876 143948 195940
rect 144012 195876 144013 195940
rect 143947 195875 144013 195876
rect 143579 188324 143645 188325
rect 143579 188260 143580 188324
rect 143644 188260 143645 188324
rect 143579 188259 143645 188260
rect 144134 186285 144194 197099
rect 144502 189005 144562 198459
rect 144499 189004 144565 189005
rect 144499 188940 144500 189004
rect 144564 188940 144565 189004
rect 144499 188939 144565 188940
rect 144131 186284 144197 186285
rect 144131 186220 144132 186284
rect 144196 186220 144197 186284
rect 144131 186219 144197 186220
rect 144686 183429 144746 199819
rect 145238 197573 145298 199819
rect 145235 197572 145301 197573
rect 145235 197508 145236 197572
rect 145300 197508 145301 197572
rect 145235 197507 145301 197508
rect 145794 183454 146414 198000
rect 146526 194610 146586 199819
rect 146891 199612 146957 199613
rect 146891 199548 146892 199612
rect 146956 199548 146957 199612
rect 146891 199547 146957 199548
rect 146526 194550 146770 194610
rect 146710 193765 146770 194550
rect 146707 193764 146773 193765
rect 146707 193700 146708 193764
rect 146772 193700 146773 193764
rect 146707 193699 146773 193700
rect 146894 186285 146954 199547
rect 147075 198388 147141 198389
rect 147075 198324 147076 198388
rect 147140 198324 147141 198388
rect 147075 198323 147141 198324
rect 147078 187509 147138 198323
rect 147446 197165 147506 199819
rect 147998 197981 148058 199819
rect 148179 199748 148245 199749
rect 148179 199684 148180 199748
rect 148244 199684 148245 199748
rect 148179 199683 148245 199684
rect 147995 197980 148061 197981
rect 147995 197916 147996 197980
rect 148060 197916 148061 197980
rect 147995 197915 148061 197916
rect 147443 197164 147509 197165
rect 147443 197100 147444 197164
rect 147508 197100 147509 197164
rect 147443 197099 147509 197100
rect 148182 190365 148242 199683
rect 148915 197980 148981 197981
rect 148915 197916 148916 197980
rect 148980 197916 148981 197980
rect 148915 197915 148981 197916
rect 148179 190364 148245 190365
rect 148179 190300 148180 190364
rect 148244 190300 148245 190364
rect 148179 190299 148245 190300
rect 148182 189141 148242 190299
rect 148179 189140 148245 189141
rect 148179 189076 148180 189140
rect 148244 189076 148245 189140
rect 148179 189075 148245 189076
rect 147075 187508 147141 187509
rect 147075 187444 147076 187508
rect 147140 187444 147141 187508
rect 147075 187443 147141 187444
rect 147078 186965 147138 187443
rect 147075 186964 147141 186965
rect 147075 186900 147076 186964
rect 147140 186900 147141 186964
rect 147075 186899 147141 186900
rect 146891 186284 146957 186285
rect 146891 186220 146892 186284
rect 146956 186220 146957 186284
rect 146891 186219 146957 186220
rect 146894 185605 146954 186219
rect 148918 185605 148978 197915
rect 149099 196756 149165 196757
rect 149099 196692 149100 196756
rect 149164 196692 149165 196756
rect 149099 196691 149165 196692
rect 149102 192949 149162 196691
rect 149470 196621 149530 199819
rect 149467 196620 149533 196621
rect 149467 196556 149468 196620
rect 149532 196556 149533 196620
rect 149467 196555 149533 196556
rect 149099 192948 149165 192949
rect 149099 192884 149100 192948
rect 149164 192884 149165 192948
rect 149099 192883 149165 192884
rect 146891 185604 146957 185605
rect 146891 185540 146892 185604
rect 146956 185540 146957 185604
rect 146891 185539 146957 185540
rect 148915 185604 148981 185605
rect 148915 185540 148916 185604
rect 148980 185540 148981 185604
rect 148915 185539 148981 185540
rect 144683 183428 144749 183429
rect 144683 183364 144684 183428
rect 144748 183364 144749 183428
rect 144683 183363 144749 183364
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141003 177988 141069 177989
rect 141003 177924 141004 177988
rect 141068 177924 141069 177988
rect 141003 177923 141069 177924
rect 137139 176356 137205 176357
rect 137139 176292 137140 176356
rect 137204 176292 137205 176356
rect 137139 176291 137205 176292
rect 135851 175948 135917 175949
rect 135851 175884 135852 175948
rect 135916 175884 135917 175948
rect 135851 175883 135917 175884
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 150022 182069 150082 199819
rect 150574 199069 150634 199819
rect 150571 199068 150637 199069
rect 150571 199004 150572 199068
rect 150636 199004 150637 199068
rect 150571 199003 150637 199004
rect 151126 198933 151186 199819
rect 151859 199748 151925 199749
rect 151859 199684 151860 199748
rect 151924 199684 151925 199748
rect 152227 199748 152293 199749
rect 152227 199746 152228 199748
rect 151859 199683 151925 199684
rect 152046 199686 152228 199746
rect 151307 199612 151373 199613
rect 151307 199548 151308 199612
rect 151372 199548 151373 199612
rect 151307 199547 151373 199548
rect 151310 198933 151370 199547
rect 151491 199068 151557 199069
rect 151491 199004 151492 199068
rect 151556 199004 151557 199068
rect 151491 199003 151557 199004
rect 151675 199068 151741 199069
rect 151675 199004 151676 199068
rect 151740 199004 151741 199068
rect 151675 199003 151741 199004
rect 151123 198932 151189 198933
rect 151123 198868 151124 198932
rect 151188 198868 151189 198932
rect 151123 198867 151189 198868
rect 151307 198932 151373 198933
rect 151307 198868 151308 198932
rect 151372 198868 151373 198932
rect 151307 198867 151373 198868
rect 150294 187954 150914 198000
rect 151123 197436 151189 197437
rect 151123 197372 151124 197436
rect 151188 197372 151189 197436
rect 151123 197371 151189 197372
rect 151126 189141 151186 197371
rect 151123 189140 151189 189141
rect 151123 189076 151124 189140
rect 151188 189076 151189 189140
rect 151123 189075 151189 189076
rect 151494 188325 151554 199003
rect 151491 188324 151557 188325
rect 151491 188260 151492 188324
rect 151556 188260 151557 188324
rect 151491 188259 151557 188260
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150019 182068 150085 182069
rect 150019 182004 150020 182068
rect 150084 182004 150085 182068
rect 150019 182003 150085 182004
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 150294 151954 150914 187398
rect 151678 181389 151738 199003
rect 151862 196757 151922 199683
rect 152046 198933 152106 199686
rect 152227 199684 152228 199686
rect 152292 199684 152293 199748
rect 152227 199683 152293 199684
rect 152043 198932 152109 198933
rect 152043 198868 152044 198932
rect 152108 198868 152109 198932
rect 152043 198867 152109 198868
rect 151859 196756 151925 196757
rect 151859 196692 151860 196756
rect 151924 196692 151925 196756
rect 151859 196691 151925 196692
rect 152598 196077 152658 200091
rect 152963 199884 153029 199885
rect 152963 199820 152964 199884
rect 153028 199820 153029 199884
rect 152963 199819 153029 199820
rect 153883 199884 153949 199885
rect 153883 199820 153884 199884
rect 153948 199820 153949 199884
rect 153883 199819 153949 199820
rect 154067 199884 154133 199885
rect 154067 199820 154068 199884
rect 154132 199820 154133 199884
rect 154067 199819 154133 199820
rect 152966 199613 153026 199819
rect 152963 199612 153029 199613
rect 152963 199548 152964 199612
rect 153028 199548 153029 199612
rect 152963 199547 153029 199548
rect 153331 199612 153397 199613
rect 153331 199548 153332 199612
rect 153396 199548 153397 199612
rect 153331 199547 153397 199548
rect 152595 196076 152661 196077
rect 152595 196012 152596 196076
rect 152660 196012 152661 196076
rect 152595 196011 152661 196012
rect 153334 191850 153394 199547
rect 153699 199204 153765 199205
rect 153699 199140 153700 199204
rect 153764 199140 153765 199204
rect 153699 199139 153765 199140
rect 153702 198750 153762 199139
rect 153886 198933 153946 199819
rect 153883 198932 153949 198933
rect 153883 198868 153884 198932
rect 153948 198868 153949 198932
rect 153883 198867 153949 198868
rect 153702 198690 153946 198750
rect 153886 196077 153946 198690
rect 154070 196213 154130 199819
rect 154254 199613 154314 200907
rect 158115 200292 158181 200293
rect 158115 200228 158116 200292
rect 158180 200228 158181 200292
rect 158115 200227 158181 200228
rect 157011 199884 157077 199885
rect 157011 199820 157012 199884
rect 157076 199820 157077 199884
rect 157011 199819 157077 199820
rect 157379 199884 157445 199885
rect 157379 199820 157380 199884
rect 157444 199820 157445 199884
rect 157379 199819 157445 199820
rect 156827 199748 156893 199749
rect 156827 199684 156828 199748
rect 156892 199684 156893 199748
rect 156827 199683 156893 199684
rect 154251 199612 154317 199613
rect 154251 199548 154252 199612
rect 154316 199548 154317 199612
rect 154251 199547 154317 199548
rect 156643 199612 156709 199613
rect 156643 199548 156644 199612
rect 156708 199548 156709 199612
rect 156643 199547 156709 199548
rect 154067 196212 154133 196213
rect 154067 196148 154068 196212
rect 154132 196148 154133 196212
rect 154067 196147 154133 196148
rect 153883 196076 153949 196077
rect 153883 196012 153884 196076
rect 153948 196012 153949 196076
rect 153883 196011 153949 196012
rect 154251 196076 154317 196077
rect 154251 196012 154252 196076
rect 154316 196012 154317 196076
rect 154251 196011 154317 196012
rect 154067 193764 154133 193765
rect 154067 193700 154068 193764
rect 154132 193700 154133 193764
rect 154067 193699 154133 193700
rect 153150 191790 153394 191850
rect 153150 191725 153210 191790
rect 153147 191724 153213 191725
rect 153147 191660 153148 191724
rect 153212 191660 153213 191724
rect 153147 191659 153213 191660
rect 154070 183157 154130 193699
rect 154067 183156 154133 183157
rect 154067 183092 154068 183156
rect 154132 183092 154133 183156
rect 154067 183091 154133 183092
rect 154254 182885 154314 196011
rect 154794 192454 155414 198000
rect 156646 196077 156706 199547
rect 156643 196076 156709 196077
rect 156643 196012 156644 196076
rect 156708 196012 156709 196076
rect 156643 196011 156709 196012
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154251 182884 154317 182885
rect 154251 182820 154252 182884
rect 154316 182820 154317 182884
rect 154251 182819 154317 182820
rect 151675 181388 151741 181389
rect 151675 181324 151676 181388
rect 151740 181324 151741 181388
rect 151675 181323 151741 181324
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 154794 156454 155414 191898
rect 156830 191181 156890 199683
rect 157014 197845 157074 199819
rect 157011 197844 157077 197845
rect 157011 197780 157012 197844
rect 157076 197780 157077 197844
rect 157011 197779 157077 197780
rect 157195 196756 157261 196757
rect 157195 196692 157196 196756
rect 157260 196692 157261 196756
rect 157195 196691 157261 196692
rect 156827 191180 156893 191181
rect 156827 191116 156828 191180
rect 156892 191116 156893 191180
rect 156827 191115 156893 191116
rect 157198 182613 157258 196691
rect 157382 196485 157442 199819
rect 158118 199749 158178 200227
rect 160326 199885 160386 201451
rect 180195 200972 180261 200973
rect 180195 200908 180196 200972
rect 180260 200908 180261 200972
rect 180195 200907 180261 200908
rect 173571 200564 173637 200565
rect 173571 200500 173572 200564
rect 173636 200500 173637 200564
rect 173571 200499 173637 200500
rect 170627 200428 170693 200429
rect 170627 200364 170628 200428
rect 170692 200364 170693 200428
rect 170627 200363 170693 200364
rect 160875 200292 160941 200293
rect 160875 200228 160876 200292
rect 160940 200228 160941 200292
rect 160875 200227 160941 200228
rect 169523 200292 169589 200293
rect 169523 200228 169524 200292
rect 169588 200228 169589 200292
rect 169523 200227 169589 200228
rect 158299 199884 158365 199885
rect 158299 199820 158300 199884
rect 158364 199820 158365 199884
rect 159403 199884 159469 199885
rect 159403 199882 159404 199884
rect 158299 199819 158365 199820
rect 159038 199822 159404 199882
rect 158115 199748 158181 199749
rect 158115 199684 158116 199748
rect 158180 199684 158181 199748
rect 158115 199683 158181 199684
rect 158302 198933 158362 199819
rect 158299 198932 158365 198933
rect 158299 198868 158300 198932
rect 158364 198868 158365 198932
rect 158299 198867 158365 198868
rect 157379 196484 157445 196485
rect 157379 196420 157380 196484
rect 157444 196420 157445 196484
rect 157379 196419 157445 196420
rect 159038 183293 159098 199822
rect 159403 199820 159404 199822
rect 159468 199820 159469 199884
rect 159403 199819 159469 199820
rect 160323 199884 160389 199885
rect 160323 199820 160324 199884
rect 160388 199820 160389 199884
rect 160323 199819 160389 199820
rect 159587 199748 159653 199749
rect 159587 199684 159588 199748
rect 159652 199684 159653 199748
rect 159587 199683 159653 199684
rect 159590 198253 159650 199683
rect 160878 199613 160938 200227
rect 163451 200156 163517 200157
rect 163451 200092 163452 200156
rect 163516 200092 163517 200156
rect 163451 200091 163517 200092
rect 163267 200020 163333 200021
rect 163267 199956 163268 200020
rect 163332 199956 163333 200020
rect 163267 199955 163333 199956
rect 161979 199884 162045 199885
rect 161979 199820 161980 199884
rect 162044 199820 162045 199884
rect 161979 199819 162045 199820
rect 160875 199612 160941 199613
rect 160875 199548 160876 199612
rect 160940 199548 160941 199612
rect 160875 199547 160941 199548
rect 161982 199341 162042 199819
rect 162531 199748 162597 199749
rect 162531 199684 162532 199748
rect 162596 199684 162597 199748
rect 162531 199683 162597 199684
rect 161979 199340 162045 199341
rect 161979 199276 161980 199340
rect 162044 199276 162045 199340
rect 161979 199275 162045 199276
rect 159587 198252 159653 198253
rect 159587 198188 159588 198252
rect 159652 198188 159653 198252
rect 159587 198187 159653 198188
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 161243 196756 161309 196757
rect 161243 196692 161244 196756
rect 161308 196692 161309 196756
rect 161243 196691 161309 196692
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159035 183292 159101 183293
rect 159035 183228 159036 183292
rect 159100 183228 159101 183292
rect 159035 183227 159101 183228
rect 157195 182612 157261 182613
rect 157195 182548 157196 182612
rect 157260 182548 157261 182612
rect 157195 182547 157261 182548
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 159294 160954 159914 196398
rect 161246 191045 161306 196691
rect 161243 191044 161309 191045
rect 161243 190980 161244 191044
rect 161308 190980 161309 191044
rect 161243 190979 161309 190980
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 161982 144261 162042 199275
rect 162534 188461 162594 199683
rect 163270 199341 163330 199955
rect 163267 199340 163333 199341
rect 163267 199276 163268 199340
rect 163332 199276 163333 199340
rect 163267 199275 163333 199276
rect 162715 198660 162781 198661
rect 162715 198596 162716 198660
rect 162780 198596 162781 198660
rect 162715 198595 162781 198596
rect 162531 188460 162597 188461
rect 162531 188396 162532 188460
rect 162596 188396 162597 188460
rect 162531 188395 162597 188396
rect 162718 184517 162778 198595
rect 163454 190093 163514 200091
rect 166579 200020 166645 200021
rect 166579 199956 166580 200020
rect 166644 199956 166645 200020
rect 166579 199955 166645 199956
rect 164003 199884 164069 199885
rect 164003 199820 164004 199884
rect 164068 199820 164069 199884
rect 164003 199819 164069 199820
rect 164555 199884 164621 199885
rect 164555 199820 164556 199884
rect 164620 199820 164621 199884
rect 164555 199819 164621 199820
rect 166395 199884 166461 199885
rect 166395 199820 166396 199884
rect 166460 199820 166461 199884
rect 166395 199819 166461 199820
rect 163635 197980 163701 197981
rect 163635 197916 163636 197980
rect 163700 197916 163701 197980
rect 163635 197915 163701 197916
rect 163451 190092 163517 190093
rect 163451 190028 163452 190092
rect 163516 190028 163517 190092
rect 163451 190027 163517 190028
rect 163638 189141 163698 197915
rect 164006 197845 164066 199819
rect 164003 197844 164069 197845
rect 164003 197780 164004 197844
rect 164068 197780 164069 197844
rect 164003 197779 164069 197780
rect 164003 197028 164069 197029
rect 164003 196964 164004 197028
rect 164068 196964 164069 197028
rect 164003 196963 164069 196964
rect 163819 196756 163885 196757
rect 163819 196692 163820 196756
rect 163884 196692 163885 196756
rect 163819 196691 163885 196692
rect 163822 190637 163882 196691
rect 163819 190636 163885 190637
rect 163819 190572 163820 190636
rect 163884 190572 163885 190636
rect 163819 190571 163885 190572
rect 163635 189140 163701 189141
rect 163635 189076 163636 189140
rect 163700 189076 163701 189140
rect 163635 189075 163701 189076
rect 162715 184516 162781 184517
rect 162715 184452 162716 184516
rect 162780 184452 162781 184516
rect 162715 184451 162781 184452
rect 164006 184381 164066 196963
rect 164371 196756 164437 196757
rect 164371 196692 164372 196756
rect 164436 196692 164437 196756
rect 164371 196691 164437 196692
rect 164374 192949 164434 196691
rect 164558 195397 164618 199819
rect 166027 199748 166093 199749
rect 166027 199684 166028 199748
rect 166092 199684 166093 199748
rect 166027 199683 166093 199684
rect 166211 199748 166277 199749
rect 166211 199684 166212 199748
rect 166276 199684 166277 199748
rect 166211 199683 166277 199684
rect 164739 199612 164805 199613
rect 164739 199548 164740 199612
rect 164804 199548 164805 199612
rect 164739 199547 164805 199548
rect 165107 199612 165173 199613
rect 165107 199548 165108 199612
rect 165172 199548 165173 199612
rect 165107 199547 165173 199548
rect 164742 198797 164802 199547
rect 164739 198796 164805 198797
rect 164739 198732 164740 198796
rect 164804 198732 164805 198796
rect 164739 198731 164805 198732
rect 164555 195396 164621 195397
rect 164555 195332 164556 195396
rect 164620 195332 164621 195396
rect 164555 195331 164621 195332
rect 164371 192948 164437 192949
rect 164371 192884 164372 192948
rect 164436 192884 164437 192948
rect 164371 192883 164437 192884
rect 164003 184380 164069 184381
rect 164003 184316 164004 184380
rect 164068 184316 164069 184380
rect 164003 184315 164069 184316
rect 165110 178669 165170 199547
rect 165475 198388 165541 198389
rect 165475 198324 165476 198388
rect 165540 198324 165541 198388
rect 165475 198323 165541 198324
rect 165478 195397 165538 198323
rect 165475 195396 165541 195397
rect 165475 195332 165476 195396
rect 165540 195332 165541 195396
rect 165475 195331 165541 195332
rect 166030 190909 166090 199683
rect 166027 190908 166093 190909
rect 166027 190844 166028 190908
rect 166092 190844 166093 190908
rect 166027 190843 166093 190844
rect 166214 178941 166274 199683
rect 166398 192541 166458 199819
rect 166395 192540 166461 192541
rect 166395 192476 166396 192540
rect 166460 192476 166461 192540
rect 166395 192475 166461 192476
rect 166582 191317 166642 199955
rect 167315 199884 167381 199885
rect 167315 199820 167316 199884
rect 167380 199820 167381 199884
rect 167315 199819 167381 199820
rect 168603 199884 168669 199885
rect 168603 199820 168604 199884
rect 168668 199820 168669 199884
rect 168603 199819 168669 199820
rect 168971 199884 169037 199885
rect 168971 199820 168972 199884
rect 169036 199820 169037 199884
rect 168971 199819 169037 199820
rect 167318 196349 167378 199819
rect 168419 199340 168485 199341
rect 168419 199276 168420 199340
rect 168484 199276 168485 199340
rect 168419 199275 168485 199276
rect 167867 198932 167933 198933
rect 167867 198868 167868 198932
rect 167932 198868 167933 198932
rect 167867 198867 167933 198868
rect 167315 196348 167381 196349
rect 167315 196284 167316 196348
rect 167380 196284 167381 196348
rect 167315 196283 167381 196284
rect 167870 191589 167930 198867
rect 168235 197708 168301 197709
rect 168235 197644 168236 197708
rect 168300 197644 168301 197708
rect 168235 197643 168301 197644
rect 167867 191588 167933 191589
rect 167867 191524 167868 191588
rect 167932 191524 167933 191588
rect 167867 191523 167933 191524
rect 166579 191316 166645 191317
rect 166579 191252 166580 191316
rect 166644 191252 166645 191316
rect 166579 191251 166645 191252
rect 168238 187101 168298 197643
rect 168422 192813 168482 199275
rect 168606 195261 168666 199819
rect 168603 195260 168669 195261
rect 168603 195196 168604 195260
rect 168668 195196 168669 195260
rect 168603 195195 168669 195196
rect 168419 192812 168485 192813
rect 168419 192748 168420 192812
rect 168484 192748 168485 192812
rect 168419 192747 168485 192748
rect 168235 187100 168301 187101
rect 168235 187036 168236 187100
rect 168300 187036 168301 187100
rect 168235 187035 168301 187036
rect 168974 184245 169034 199819
rect 169339 199748 169405 199749
rect 169339 199684 169340 199748
rect 169404 199684 169405 199748
rect 169339 199683 169405 199684
rect 169155 199612 169221 199613
rect 169155 199548 169156 199612
rect 169220 199548 169221 199612
rect 169155 199547 169221 199548
rect 169158 186013 169218 199547
rect 169342 186829 169402 199683
rect 169526 199613 169586 200227
rect 170630 199885 170690 200363
rect 170995 200156 171061 200157
rect 170995 200092 170996 200156
rect 171060 200092 171061 200156
rect 170995 200091 171061 200092
rect 170627 199884 170693 199885
rect 170627 199820 170628 199884
rect 170692 199820 170693 199884
rect 170627 199819 170693 199820
rect 169523 199612 169589 199613
rect 169523 199548 169524 199612
rect 169588 199548 169589 199612
rect 169523 199547 169589 199548
rect 170811 199612 170877 199613
rect 170811 199548 170812 199612
rect 170876 199548 170877 199612
rect 170811 199547 170877 199548
rect 169707 197572 169773 197573
rect 169707 197508 169708 197572
rect 169772 197508 169773 197572
rect 169707 197507 169773 197508
rect 169710 187645 169770 197507
rect 170814 197437 170874 199547
rect 170811 197436 170877 197437
rect 170811 197372 170812 197436
rect 170876 197372 170877 197436
rect 170811 197371 170877 197372
rect 170998 196757 171058 200091
rect 173203 200020 173269 200021
rect 173203 199956 173204 200020
rect 173268 199956 173269 200020
rect 173203 199955 173269 199956
rect 171363 199884 171429 199885
rect 171363 199820 171364 199884
rect 171428 199820 171429 199884
rect 171363 199819 171429 199820
rect 172283 199884 172349 199885
rect 172283 199820 172284 199884
rect 172348 199820 172349 199884
rect 172283 199819 172349 199820
rect 171366 197573 171426 199819
rect 171363 197572 171429 197573
rect 171363 197508 171364 197572
rect 171428 197508 171429 197572
rect 171363 197507 171429 197508
rect 170995 196756 171061 196757
rect 170995 196692 170996 196756
rect 171060 196692 171061 196756
rect 170995 196691 171061 196692
rect 171731 196484 171797 196485
rect 171731 196420 171732 196484
rect 171796 196420 171797 196484
rect 171731 196419 171797 196420
rect 169707 187644 169773 187645
rect 169707 187580 169708 187644
rect 169772 187580 169773 187644
rect 169707 187579 169773 187580
rect 169339 186828 169405 186829
rect 169339 186764 169340 186828
rect 169404 186764 169405 186828
rect 169339 186763 169405 186764
rect 169155 186012 169221 186013
rect 169155 185948 169156 186012
rect 169220 185948 169221 186012
rect 169155 185947 169221 185948
rect 168971 184244 169037 184245
rect 168971 184180 168972 184244
rect 169036 184180 169037 184244
rect 168971 184179 169037 184180
rect 166211 178940 166277 178941
rect 166211 178876 166212 178940
rect 166276 178876 166277 178940
rect 166211 178875 166277 178876
rect 171734 178805 171794 196419
rect 172286 189821 172346 199819
rect 173206 193230 173266 199955
rect 173574 198933 173634 200499
rect 180198 200021 180258 200907
rect 180195 200020 180261 200021
rect 180195 199956 180196 200020
rect 180260 199956 180261 200020
rect 180195 199955 180261 199956
rect 174307 199884 174373 199885
rect 174307 199820 174308 199884
rect 174372 199820 174373 199884
rect 174307 199819 174373 199820
rect 174675 199884 174741 199885
rect 174675 199820 174676 199884
rect 174740 199820 174741 199884
rect 174675 199819 174741 199820
rect 176331 199884 176397 199885
rect 176331 199820 176332 199884
rect 176396 199820 176397 199884
rect 176331 199819 176397 199820
rect 173571 198932 173637 198933
rect 173571 198868 173572 198932
rect 173636 198868 173637 198932
rect 173571 198867 173637 198868
rect 173387 198660 173453 198661
rect 173387 198596 173388 198660
rect 173452 198596 173453 198660
rect 173387 198595 173453 198596
rect 173755 198660 173821 198661
rect 173755 198596 173756 198660
rect 173820 198596 173821 198660
rect 173755 198595 173821 198596
rect 173390 197029 173450 198595
rect 173387 197028 173453 197029
rect 173387 196964 173388 197028
rect 173452 196964 173453 197028
rect 173387 196963 173453 196964
rect 173022 193170 173266 193230
rect 173022 193085 173082 193170
rect 173019 193084 173085 193085
rect 173019 193020 173020 193084
rect 173084 193020 173085 193084
rect 173019 193019 173085 193020
rect 172283 189820 172349 189821
rect 172283 189756 172284 189820
rect 172348 189756 172349 189820
rect 172283 189755 172349 189756
rect 173758 185877 173818 198595
rect 174310 197370 174370 199819
rect 174678 198661 174738 199819
rect 176334 199477 176394 199819
rect 175411 199476 175477 199477
rect 175411 199412 175412 199476
rect 175476 199412 175477 199476
rect 175411 199411 175477 199412
rect 176331 199476 176397 199477
rect 176331 199412 176332 199476
rect 176396 199412 176397 199476
rect 176331 199411 176397 199412
rect 174675 198660 174741 198661
rect 174675 198596 174676 198660
rect 174740 198596 174741 198660
rect 174675 198595 174741 198596
rect 174310 197310 174554 197370
rect 173755 185876 173821 185877
rect 173755 185812 173756 185876
rect 173820 185812 173821 185876
rect 173755 185811 173821 185812
rect 174494 185741 174554 197310
rect 174675 196076 174741 196077
rect 174675 196012 174676 196076
rect 174740 196012 174741 196076
rect 174675 196011 174741 196012
rect 174678 187373 174738 196011
rect 174859 195804 174925 195805
rect 174859 195740 174860 195804
rect 174924 195740 174925 195804
rect 174859 195739 174925 195740
rect 174675 187372 174741 187373
rect 174675 187308 174676 187372
rect 174740 187308 174741 187372
rect 174675 187307 174741 187308
rect 174862 187237 174922 195739
rect 175227 193220 175293 193221
rect 175227 193156 175228 193220
rect 175292 193156 175293 193220
rect 175227 193155 175293 193156
rect 174859 187236 174925 187237
rect 174859 187172 174860 187236
rect 174924 187172 174925 187236
rect 174859 187171 174925 187172
rect 175230 186149 175290 193155
rect 175414 190229 175474 199411
rect 176515 197436 176581 197437
rect 176515 197372 176516 197436
rect 176580 197372 176581 197436
rect 176515 197371 176581 197372
rect 175411 190228 175477 190229
rect 175411 190164 175412 190228
rect 175476 190164 175477 190228
rect 175411 190163 175477 190164
rect 175414 189141 175474 190163
rect 175411 189140 175477 189141
rect 175411 189076 175412 189140
rect 175476 189076 175477 189140
rect 175411 189075 175477 189076
rect 176518 188597 176578 197371
rect 176515 188596 176581 188597
rect 176515 188532 176516 188596
rect 176580 188532 176581 188596
rect 176515 188531 176581 188532
rect 175227 186148 175293 186149
rect 175227 186084 175228 186148
rect 175292 186084 175293 186148
rect 175227 186083 175293 186084
rect 174491 185740 174557 185741
rect 174491 185676 174492 185740
rect 174556 185676 174557 185740
rect 174491 185675 174557 185676
rect 177294 178954 177914 198000
rect 171731 178804 171797 178805
rect 171731 178740 171732 178804
rect 171796 178740 171797 178804
rect 171731 178739 171797 178740
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 165107 178668 165173 178669
rect 165107 178604 165108 178668
rect 165172 178604 165173 178668
rect 165107 178603 165173 178604
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 161979 144260 162045 144261
rect 161979 144196 161980 144260
rect 162044 144196 162045 144260
rect 161979 144195 162045 144196
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181486 141405 181546 201723
rect 184979 201516 185045 201517
rect 184979 201452 184980 201516
rect 185044 201452 185045 201516
rect 184979 201451 185045 201452
rect 184982 199205 185042 201451
rect 186822 200973 186882 233275
rect 186819 200972 186885 200973
rect 186819 200908 186820 200972
rect 186884 200908 186885 200972
rect 186819 200907 186885 200908
rect 184979 199204 185045 199205
rect 184979 199140 184980 199204
rect 185044 199140 185045 199204
rect 184979 199139 185045 199140
rect 181794 183454 182414 198000
rect 185347 197980 185413 197981
rect 185347 197916 185348 197980
rect 185412 197916 185413 197980
rect 185347 197915 185413 197916
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 181483 141404 181549 141405
rect 181483 141340 181484 141404
rect 181548 141340 181549 141404
rect 181483 141339 181549 141340
rect 134379 140316 134445 140317
rect 134379 140252 134380 140316
rect 134444 140252 134445 140316
rect 134379 140251 134445 140252
rect 126099 139364 126165 139365
rect 126099 139300 126100 139364
rect 126164 139300 126165 139364
rect 126099 139299 126165 139300
rect 136955 139364 137021 139365
rect 136955 139300 136956 139364
rect 137020 139300 137021 139364
rect 136955 139299 137021 139300
rect 126102 138549 126162 139299
rect 136958 138821 137018 139299
rect 136955 138820 137021 138821
rect 136955 138756 136956 138820
rect 137020 138756 137021 138820
rect 136955 138755 137021 138756
rect 126099 138548 126165 138549
rect 126099 138484 126100 138548
rect 126164 138484 126165 138548
rect 126099 138483 126165 138484
rect 185350 138277 185410 197915
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 185715 183020 185781 183021
rect 185715 182956 185716 183020
rect 185780 182956 185781 183020
rect 185715 182955 185781 182956
rect 185347 138276 185413 138277
rect 185347 138212 185348 138276
rect 185412 138212 185413 138276
rect 185347 138211 185413 138212
rect 185718 137869 185778 182955
rect 186083 182884 186149 182885
rect 186083 182820 186084 182884
rect 186148 182820 186149 182884
rect 186083 182819 186149 182820
rect 124811 137868 124877 137869
rect 124811 137804 124812 137868
rect 124876 137804 124877 137868
rect 124811 137803 124877 137804
rect 185715 137868 185781 137869
rect 185715 137804 185716 137868
rect 185780 137804 185781 137868
rect 185715 137803 185781 137804
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 186086 91221 186146 182819
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 187006 143173 187066 259251
rect 187190 143445 187250 259931
rect 188291 245716 188357 245717
rect 188291 245652 188292 245716
rect 188356 245652 188357 245716
rect 188291 245651 188357 245652
rect 188294 200837 188354 245651
rect 188475 218108 188541 218109
rect 188475 218044 188476 218108
rect 188540 218044 188541 218108
rect 188475 218043 188541 218044
rect 188291 200836 188357 200837
rect 188291 200772 188292 200836
rect 188356 200772 188357 200836
rect 188291 200771 188357 200772
rect 188478 199749 188538 218043
rect 188475 199748 188541 199749
rect 188475 199684 188476 199748
rect 188540 199684 188541 199748
rect 188475 199683 188541 199684
rect 190499 196620 190565 196621
rect 190499 196556 190500 196620
rect 190564 196556 190565 196620
rect 190499 196555 190565 196556
rect 189027 190772 189093 190773
rect 189027 190708 189028 190772
rect 189092 190708 189093 190772
rect 189027 190707 189093 190708
rect 187739 189956 187805 189957
rect 187739 189892 187740 189956
rect 187804 189892 187805 189956
rect 187739 189891 187805 189892
rect 187742 189685 187802 189891
rect 187739 189684 187805 189685
rect 187739 189620 187740 189684
rect 187804 189620 187805 189684
rect 187739 189619 187805 189620
rect 187187 143444 187253 143445
rect 187187 143380 187188 143444
rect 187252 143380 187253 143444
rect 187187 143379 187253 143380
rect 187003 143172 187069 143173
rect 187003 143108 187004 143172
rect 187068 143108 187069 143172
rect 187003 143107 187069 143108
rect 187371 140180 187437 140181
rect 187371 140116 187372 140180
rect 187436 140116 187437 140180
rect 187371 140115 187437 140116
rect 187187 139364 187253 139365
rect 187187 139300 187188 139364
rect 187252 139300 187253 139364
rect 187187 139299 187253 139300
rect 187003 139228 187069 139229
rect 187003 139164 187004 139228
rect 187068 139164 187069 139228
rect 187003 139163 187069 139164
rect 186267 138276 186333 138277
rect 186267 138212 186268 138276
rect 186332 138212 186333 138276
rect 186267 138211 186333 138212
rect 186270 134469 186330 138211
rect 186819 136644 186885 136645
rect 186819 136580 186820 136644
rect 186884 136580 186885 136644
rect 186819 136579 186885 136580
rect 186267 134468 186333 134469
rect 186267 134404 186268 134468
rect 186332 134404 186333 134468
rect 186267 134403 186333 134404
rect 186083 91220 186149 91221
rect 186083 91156 186084 91220
rect 186148 91156 186149 91220
rect 186083 91155 186149 91156
rect 186083 82244 186149 82245
rect 186083 82180 186084 82244
rect 186148 82180 186149 82244
rect 186083 82179 186149 82180
rect 135851 81972 135917 81973
rect 135851 81908 135852 81972
rect 135916 81908 135917 81972
rect 135851 81907 135917 81908
rect 176699 81972 176765 81973
rect 176699 81908 176700 81972
rect 176764 81908 176765 81972
rect 176699 81907 176765 81908
rect 131435 81292 131501 81293
rect 131435 81228 131436 81292
rect 131500 81228 131501 81292
rect 131435 81227 131501 81228
rect 131438 80069 131498 81227
rect 133275 81156 133341 81157
rect 133275 81092 133276 81156
rect 133340 81092 133341 81156
rect 133275 81091 133341 81092
rect 131435 80068 131501 80069
rect 131435 80004 131436 80068
rect 131500 80004 131501 80068
rect 131435 80003 131501 80004
rect 133278 79933 133338 81091
rect 135483 81020 135549 81021
rect 135483 80956 135484 81020
rect 135548 80956 135549 81020
rect 135483 80955 135549 80956
rect 134379 80748 134445 80749
rect 134379 80684 134380 80748
rect 134444 80684 134445 80748
rect 134379 80683 134445 80684
rect 134382 79933 134442 80683
rect 133275 79932 133341 79933
rect 133275 79868 133276 79932
rect 133340 79868 133341 79932
rect 133275 79867 133341 79868
rect 134379 79932 134445 79933
rect 134379 79868 134380 79932
rect 134444 79868 134445 79932
rect 134379 79867 134445 79868
rect 135115 79932 135181 79933
rect 135115 79868 135116 79932
rect 135180 79868 135181 79932
rect 135115 79867 135181 79868
rect 134931 79796 134997 79797
rect 134931 79732 134932 79796
rect 134996 79732 134997 79796
rect 134931 79731 134997 79732
rect 134934 78573 134994 79731
rect 135118 79117 135178 79867
rect 135299 79796 135365 79797
rect 135299 79732 135300 79796
rect 135364 79732 135365 79796
rect 135299 79731 135365 79732
rect 135115 79116 135181 79117
rect 135115 79052 135116 79116
rect 135180 79052 135181 79116
rect 135115 79051 135181 79052
rect 134931 78572 134997 78573
rect 134931 78508 134932 78572
rect 134996 78508 134997 78572
rect 134931 78507 134997 78508
rect 124075 78164 124141 78165
rect 124075 78100 124076 78164
rect 124140 78100 124141 78164
rect 124075 78099 124141 78100
rect 122971 67012 123037 67013
rect 122971 66948 122972 67012
rect 123036 66948 123037 67012
rect 122971 66947 123037 66948
rect 122051 64292 122117 64293
rect 122051 64228 122052 64292
rect 122116 64228 122117 64292
rect 122051 64227 122117 64228
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133091 75988 133157 75989
rect 133091 75924 133092 75988
rect 133156 75924 133157 75988
rect 133091 75923 133157 75924
rect 133094 70957 133154 75923
rect 133091 70956 133157 70957
rect 133091 70892 133092 70956
rect 133156 70892 133157 70956
rect 133091 70891 133157 70892
rect 135302 69869 135362 79731
rect 135486 79117 135546 80955
rect 135667 79932 135733 79933
rect 135667 79868 135668 79932
rect 135732 79868 135733 79932
rect 135667 79867 135733 79868
rect 135483 79116 135549 79117
rect 135483 79052 135484 79116
rect 135548 79052 135549 79116
rect 135483 79051 135549 79052
rect 135670 78437 135730 79867
rect 135854 79797 135914 81907
rect 137323 81836 137389 81837
rect 137323 81772 137324 81836
rect 137388 81772 137389 81836
rect 137323 81771 137389 81772
rect 175043 81836 175109 81837
rect 175043 81772 175044 81836
rect 175108 81772 175109 81836
rect 175043 81771 175109 81772
rect 137326 79933 137386 81771
rect 141371 81428 141437 81429
rect 141371 81364 141372 81428
rect 141436 81364 141437 81428
rect 141371 81363 141437 81364
rect 136403 79932 136469 79933
rect 136403 79868 136404 79932
rect 136468 79868 136469 79932
rect 136403 79867 136469 79868
rect 137323 79932 137389 79933
rect 137323 79868 137324 79932
rect 137388 79868 137389 79932
rect 137323 79867 137389 79868
rect 138611 79932 138677 79933
rect 138611 79868 138612 79932
rect 138676 79868 138677 79932
rect 138611 79867 138677 79868
rect 140083 79932 140149 79933
rect 140083 79868 140084 79932
rect 140148 79868 140149 79932
rect 140083 79867 140149 79868
rect 140267 79932 140333 79933
rect 140267 79868 140268 79932
rect 140332 79868 140333 79932
rect 140267 79867 140333 79868
rect 141187 79932 141253 79933
rect 141187 79868 141188 79932
rect 141252 79868 141253 79932
rect 141187 79867 141253 79868
rect 135851 79796 135917 79797
rect 135851 79732 135852 79796
rect 135916 79732 135917 79796
rect 135851 79731 135917 79732
rect 136219 79796 136285 79797
rect 136219 79732 136220 79796
rect 136284 79732 136285 79796
rect 136219 79731 136285 79732
rect 135667 78436 135733 78437
rect 135667 78372 135668 78436
rect 135732 78372 135733 78436
rect 135667 78371 135733 78372
rect 135851 77756 135917 77757
rect 135851 77692 135852 77756
rect 135916 77692 135917 77756
rect 135851 77691 135917 77692
rect 135299 69868 135365 69869
rect 135299 69804 135300 69868
rect 135364 69804 135365 69868
rect 135299 69803 135365 69804
rect 135854 67149 135914 77691
rect 136222 76125 136282 79731
rect 136219 76124 136285 76125
rect 136219 76060 136220 76124
rect 136284 76060 136285 76124
rect 136219 76059 136285 76060
rect 136406 75989 136466 79867
rect 138059 79524 138125 79525
rect 138059 79460 138060 79524
rect 138124 79460 138125 79524
rect 138059 79459 138125 79460
rect 136771 79116 136837 79117
rect 136771 79052 136772 79116
rect 136836 79052 136837 79116
rect 136771 79051 136837 79052
rect 136774 78690 136834 79051
rect 136590 78630 136834 78690
rect 136403 75988 136469 75989
rect 136403 75924 136404 75988
rect 136468 75924 136469 75988
rect 136403 75923 136469 75924
rect 136590 71365 136650 78630
rect 136587 71364 136653 71365
rect 136587 71300 136588 71364
rect 136652 71300 136653 71364
rect 136587 71299 136653 71300
rect 135851 67148 135917 67149
rect 135851 67084 135852 67148
rect 135916 67084 135917 67148
rect 135851 67083 135917 67084
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 138062 65925 138122 79459
rect 138614 79389 138674 79867
rect 139347 79796 139413 79797
rect 139347 79732 139348 79796
rect 139412 79732 139413 79796
rect 139347 79731 139413 79732
rect 138611 79388 138677 79389
rect 138611 79324 138612 79388
rect 138676 79324 138677 79388
rect 138611 79323 138677 79324
rect 139350 79253 139410 79731
rect 139347 79252 139413 79253
rect 139347 79188 139348 79252
rect 139412 79188 139413 79252
rect 139347 79187 139413 79188
rect 139899 79116 139965 79117
rect 139899 79052 139900 79116
rect 139964 79052 139965 79116
rect 139899 79051 139965 79052
rect 139347 78028 139413 78029
rect 139347 77964 139348 78028
rect 139412 77964 139413 78028
rect 139347 77963 139413 77964
rect 138243 77620 138309 77621
rect 138243 77556 138244 77620
rect 138308 77556 138309 77620
rect 138243 77555 138309 77556
rect 138246 67421 138306 77555
rect 139350 72317 139410 77963
rect 139347 72316 139413 72317
rect 139347 72252 139348 72316
rect 139412 72252 139413 72316
rect 139347 72251 139413 72252
rect 139902 69597 139962 79051
rect 140086 76397 140146 79867
rect 140270 76805 140330 79867
rect 140635 79796 140701 79797
rect 140635 79732 140636 79796
rect 140700 79732 140701 79796
rect 140635 79731 140701 79732
rect 140451 78572 140517 78573
rect 140451 78508 140452 78572
rect 140516 78508 140517 78572
rect 140451 78507 140517 78508
rect 140267 76804 140333 76805
rect 140267 76740 140268 76804
rect 140332 76740 140333 76804
rect 140267 76739 140333 76740
rect 140083 76396 140149 76397
rect 140083 76332 140084 76396
rect 140148 76332 140149 76396
rect 140083 76331 140149 76332
rect 140454 73949 140514 78507
rect 140638 75445 140698 79731
rect 141190 78165 141250 79867
rect 141374 79661 141434 81363
rect 166579 81292 166645 81293
rect 166579 81228 166580 81292
rect 166644 81228 166645 81292
rect 166579 81227 166645 81228
rect 147443 80884 147509 80885
rect 147443 80820 147444 80884
rect 147508 80820 147509 80884
rect 147443 80819 147509 80820
rect 154803 80884 154869 80885
rect 154803 80820 154804 80884
rect 154868 80820 154869 80884
rect 154803 80819 154869 80820
rect 147446 79933 147506 80819
rect 154251 80204 154317 80205
rect 154251 80140 154252 80204
rect 154316 80140 154317 80204
rect 154251 80139 154317 80140
rect 144499 79932 144565 79933
rect 144499 79868 144500 79932
rect 144564 79868 144565 79932
rect 144499 79867 144565 79868
rect 147443 79932 147509 79933
rect 147443 79868 147444 79932
rect 147508 79868 147509 79932
rect 147443 79867 147509 79868
rect 148547 79932 148613 79933
rect 148547 79868 148548 79932
rect 148612 79868 148613 79932
rect 149467 79932 149533 79933
rect 149467 79930 149468 79932
rect 148547 79867 148613 79868
rect 149286 79870 149468 79930
rect 141371 79660 141437 79661
rect 141371 79596 141372 79660
rect 141436 79596 141437 79660
rect 141371 79595 141437 79596
rect 143947 79660 144013 79661
rect 143947 79596 143948 79660
rect 144012 79596 144013 79660
rect 143947 79595 144013 79596
rect 142659 79116 142725 79117
rect 142659 79052 142660 79116
rect 142724 79052 142725 79116
rect 142659 79051 142725 79052
rect 142107 78436 142173 78437
rect 142107 78372 142108 78436
rect 142172 78372 142173 78436
rect 142107 78371 142173 78372
rect 141187 78164 141253 78165
rect 141187 78100 141188 78164
rect 141252 78100 141253 78164
rect 141187 78099 141253 78100
rect 140635 75444 140701 75445
rect 140635 75380 140636 75444
rect 140700 75380 140701 75444
rect 140635 75379 140701 75380
rect 140451 73948 140517 73949
rect 140451 73884 140452 73948
rect 140516 73884 140517 73948
rect 140451 73883 140517 73884
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 142110 70413 142170 78371
rect 142662 72861 142722 79051
rect 143579 77892 143645 77893
rect 143579 77828 143580 77892
rect 143644 77828 143645 77892
rect 143579 77827 143645 77828
rect 142659 72860 142725 72861
rect 142659 72796 142660 72860
rect 142724 72796 142725 72860
rect 142659 72795 142725 72796
rect 139899 69596 139965 69597
rect 139899 69532 139900 69596
rect 139964 69532 139965 69596
rect 139899 69531 139965 69532
rect 138243 67420 138309 67421
rect 138243 67356 138244 67420
rect 138308 67356 138309 67420
rect 138243 67355 138309 67356
rect 134931 63884 134997 63885
rect 134931 63820 134932 63884
rect 134996 63820 134997 63884
rect 134931 63819 134997 63820
rect 134934 62117 134994 63819
rect 134931 62116 134997 62117
rect 134931 62052 134932 62116
rect 134996 62052 134997 62116
rect 134931 62051 134997 62052
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 138059 65924 138125 65925
rect 138059 65860 138060 65924
rect 138124 65860 138125 65924
rect 138059 65859 138125 65860
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 142107 70412 142173 70413
rect 142107 70348 142108 70412
rect 142172 70348 142173 70412
rect 142107 70347 142173 70348
rect 143582 68509 143642 77827
rect 143950 75717 144010 79595
rect 144502 78165 144562 79867
rect 145051 79660 145117 79661
rect 145051 79596 145052 79660
rect 145116 79596 145117 79660
rect 145051 79595 145117 79596
rect 144499 78164 144565 78165
rect 144499 78100 144500 78164
rect 144564 78100 144565 78164
rect 144499 78099 144565 78100
rect 144131 77756 144197 77757
rect 144131 77692 144132 77756
rect 144196 77692 144197 77756
rect 144131 77691 144197 77692
rect 143947 75716 144013 75717
rect 143947 75652 143948 75716
rect 144012 75652 144013 75716
rect 143947 75651 144013 75652
rect 143579 68508 143645 68509
rect 143579 68444 143580 68508
rect 143644 68444 143645 68508
rect 143579 68443 143645 68444
rect 144134 64837 144194 77691
rect 145054 69733 145114 79595
rect 147811 79388 147877 79389
rect 147811 79324 147812 79388
rect 147876 79324 147877 79388
rect 147811 79323 147877 79324
rect 146707 78028 146773 78029
rect 145794 75454 146414 78000
rect 146707 77964 146708 78028
rect 146772 77964 146773 78028
rect 146707 77963 146773 77964
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 146710 75309 146770 77963
rect 146707 75308 146773 75309
rect 146707 75244 146708 75308
rect 146772 75244 146773 75308
rect 146707 75243 146773 75244
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145051 69732 145117 69733
rect 145051 69668 145052 69732
rect 145116 69668 145117 69732
rect 145051 69667 145117 69668
rect 144131 64836 144197 64837
rect 144131 64772 144132 64836
rect 144196 64772 144197 64836
rect 144131 64771 144197 64772
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 39454 146414 74898
rect 147814 64429 147874 79323
rect 147995 78300 148061 78301
rect 147995 78236 147996 78300
rect 148060 78236 148061 78300
rect 147995 78235 148061 78236
rect 147811 64428 147877 64429
rect 147811 64364 147812 64428
rect 147876 64364 147877 64428
rect 147811 64363 147877 64364
rect 147998 64293 148058 78235
rect 148550 76261 148610 79867
rect 149286 78437 149346 79870
rect 149467 79868 149468 79870
rect 149532 79868 149533 79932
rect 149467 79867 149533 79868
rect 150939 79932 151005 79933
rect 150939 79868 150940 79932
rect 151004 79868 151005 79932
rect 150939 79867 151005 79868
rect 152595 79932 152661 79933
rect 152595 79868 152596 79932
rect 152660 79868 152661 79932
rect 152595 79867 152661 79868
rect 152779 79932 152845 79933
rect 152779 79868 152780 79932
rect 152844 79868 152845 79932
rect 152779 79867 152845 79868
rect 153699 79932 153765 79933
rect 153699 79868 153700 79932
rect 153764 79868 153765 79932
rect 153699 79867 153765 79868
rect 154067 79932 154133 79933
rect 154067 79868 154068 79932
rect 154132 79868 154133 79932
rect 154254 79930 154314 80139
rect 154254 79870 154498 79930
rect 154067 79867 154133 79868
rect 149283 78436 149349 78437
rect 149283 78372 149284 78436
rect 149348 78372 149349 78436
rect 149283 78371 149349 78372
rect 150942 78301 151002 79867
rect 151123 79796 151189 79797
rect 151123 79732 151124 79796
rect 151188 79732 151189 79796
rect 151123 79731 151189 79732
rect 150939 78300 151005 78301
rect 150939 78236 150940 78300
rect 151004 78236 151005 78300
rect 150939 78235 151005 78236
rect 149283 78028 149349 78029
rect 149283 77964 149284 78028
rect 149348 77964 149349 78028
rect 149283 77963 149349 77964
rect 149651 78028 149717 78029
rect 149651 77964 149652 78028
rect 149716 77964 149717 78028
rect 149651 77963 149717 77964
rect 148547 76260 148613 76261
rect 148547 76196 148548 76260
rect 148612 76196 148613 76260
rect 148547 76195 148613 76196
rect 149286 71229 149346 77963
rect 149654 71773 149714 77963
rect 149651 71772 149717 71773
rect 149651 71708 149652 71772
rect 149716 71708 149717 71772
rect 149651 71707 149717 71708
rect 149283 71228 149349 71229
rect 149283 71164 149284 71228
rect 149348 71164 149349 71228
rect 149283 71163 149349 71164
rect 147995 64292 148061 64293
rect 147995 64228 147996 64292
rect 148060 64228 148061 64292
rect 147995 64227 148061 64228
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 78000
rect 151126 73133 151186 79731
rect 152598 74357 152658 79867
rect 152782 77893 152842 79867
rect 153702 78029 153762 79867
rect 154070 78709 154130 79867
rect 154251 79796 154317 79797
rect 154251 79732 154252 79796
rect 154316 79732 154317 79796
rect 154251 79731 154317 79732
rect 154067 78708 154133 78709
rect 154067 78644 154068 78708
rect 154132 78644 154133 78708
rect 154067 78643 154133 78644
rect 153699 78028 153765 78029
rect 153699 77964 153700 78028
rect 153764 77964 153765 78028
rect 153699 77963 153765 77964
rect 152779 77892 152845 77893
rect 152779 77828 152780 77892
rect 152844 77828 152845 77892
rect 152779 77827 152845 77828
rect 152595 74356 152661 74357
rect 152595 74292 152596 74356
rect 152660 74292 152661 74356
rect 152595 74291 152661 74292
rect 151123 73132 151189 73133
rect 151123 73068 151124 73132
rect 151188 73068 151189 73132
rect 151123 73067 151189 73068
rect 154254 69869 154314 79731
rect 154251 69868 154317 69869
rect 154251 69804 154252 69868
rect 154316 69804 154317 69868
rect 154251 69803 154317 69804
rect 154438 65381 154498 79870
rect 154806 79661 154866 80819
rect 161059 80204 161125 80205
rect 161059 80140 161060 80204
rect 161124 80140 161125 80204
rect 161059 80139 161125 80140
rect 160507 79932 160573 79933
rect 160507 79868 160508 79932
rect 160572 79868 160573 79932
rect 160507 79867 160573 79868
rect 158483 79796 158549 79797
rect 158483 79732 158484 79796
rect 158548 79732 158549 79796
rect 158483 79731 158549 79732
rect 158851 79796 158917 79797
rect 158851 79732 158852 79796
rect 158916 79732 158917 79796
rect 158851 79731 158917 79732
rect 159587 79796 159653 79797
rect 159587 79732 159588 79796
rect 159652 79732 159653 79796
rect 159587 79731 159653 79732
rect 154803 79660 154869 79661
rect 154803 79596 154804 79660
rect 154868 79596 154869 79660
rect 154803 79595 154869 79596
rect 156091 78708 156157 78709
rect 156091 78644 156092 78708
rect 156156 78644 156157 78708
rect 156091 78643 156157 78644
rect 154435 65380 154501 65381
rect 154435 65316 154436 65380
rect 154500 65316 154501 65380
rect 154435 65315 154501 65316
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 78000
rect 156094 74221 156154 78643
rect 156643 78572 156709 78573
rect 156643 78508 156644 78572
rect 156708 78508 156709 78572
rect 156643 78507 156709 78508
rect 156091 74220 156157 74221
rect 156091 74156 156092 74220
rect 156156 74156 156157 74220
rect 156091 74155 156157 74156
rect 156646 73133 156706 78507
rect 158115 76668 158181 76669
rect 158115 76604 158116 76668
rect 158180 76604 158181 76668
rect 158115 76603 158181 76604
rect 158299 76668 158365 76669
rect 158299 76604 158300 76668
rect 158364 76604 158365 76668
rect 158299 76603 158365 76604
rect 156643 73132 156709 73133
rect 156643 73068 156644 73132
rect 156708 73068 156709 73132
rect 156643 73067 156709 73068
rect 158118 65925 158178 76603
rect 158302 69597 158362 76603
rect 158486 72725 158546 79731
rect 158854 75989 158914 79731
rect 159590 78573 159650 79731
rect 159587 78572 159653 78573
rect 159587 78508 159588 78572
rect 159652 78508 159653 78572
rect 159587 78507 159653 78508
rect 158851 75988 158917 75989
rect 158851 75924 158852 75988
rect 158916 75924 158917 75988
rect 158851 75923 158917 75924
rect 158483 72724 158549 72725
rect 158483 72660 158484 72724
rect 158548 72660 158549 72724
rect 158483 72659 158549 72660
rect 158299 69596 158365 69597
rect 158299 69532 158300 69596
rect 158364 69532 158365 69596
rect 158299 69531 158365 69532
rect 158115 65924 158181 65925
rect 158115 65860 158116 65924
rect 158180 65860 158181 65924
rect 158115 65859 158181 65860
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 78000
rect 160510 75989 160570 79867
rect 160691 77212 160757 77213
rect 160691 77148 160692 77212
rect 160756 77148 160757 77212
rect 160691 77147 160757 77148
rect 160507 75988 160573 75989
rect 160507 75924 160508 75988
rect 160572 75924 160573 75988
rect 160507 75923 160573 75924
rect 160694 66061 160754 77147
rect 161062 66197 161122 80139
rect 161795 79932 161861 79933
rect 161795 79868 161796 79932
rect 161860 79868 161861 79932
rect 161795 79867 161861 79868
rect 162347 79932 162413 79933
rect 162347 79868 162348 79932
rect 162412 79868 162413 79932
rect 162347 79867 162413 79868
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 161243 78708 161309 78709
rect 161243 78644 161244 78708
rect 161308 78644 161309 78708
rect 161243 78643 161309 78644
rect 161059 66196 161125 66197
rect 161059 66132 161060 66196
rect 161124 66132 161125 66196
rect 161059 66131 161125 66132
rect 160691 66060 160757 66061
rect 160691 65996 160692 66060
rect 160756 65996 160757 66060
rect 160691 65995 160757 65996
rect 161246 63477 161306 78643
rect 161798 73677 161858 79867
rect 161979 78164 162045 78165
rect 161979 78100 161980 78164
rect 162044 78100 162045 78164
rect 161979 78099 162045 78100
rect 161795 73676 161861 73677
rect 161795 73612 161796 73676
rect 161860 73612 161861 73676
rect 161795 73611 161861 73612
rect 161982 65789 162042 78099
rect 162350 74493 162410 79867
rect 162715 79524 162781 79525
rect 162715 79460 162716 79524
rect 162780 79460 162781 79524
rect 162715 79459 162781 79460
rect 162347 74492 162413 74493
rect 162347 74428 162348 74492
rect 162412 74428 162413 74492
rect 162347 74427 162413 74428
rect 162718 67013 162778 79459
rect 163454 78709 163514 79867
rect 163635 79796 163701 79797
rect 163635 79732 163636 79796
rect 163700 79732 163701 79796
rect 163635 79731 163701 79732
rect 164555 79796 164621 79797
rect 164555 79732 164556 79796
rect 164620 79732 164621 79796
rect 164555 79731 164621 79732
rect 163451 78708 163517 78709
rect 163451 78644 163452 78708
rect 163516 78644 163517 78708
rect 163451 78643 163517 78644
rect 162899 77620 162965 77621
rect 162899 77556 162900 77620
rect 162964 77556 162965 77620
rect 162899 77555 162965 77556
rect 162902 70957 162962 77555
rect 163451 75852 163517 75853
rect 163451 75788 163452 75852
rect 163516 75788 163517 75852
rect 163451 75787 163517 75788
rect 162899 70956 162965 70957
rect 162899 70892 162900 70956
rect 162964 70892 162965 70956
rect 162899 70891 162965 70892
rect 162715 67012 162781 67013
rect 162715 66948 162716 67012
rect 162780 66948 162781 67012
rect 162715 66947 162781 66948
rect 161979 65788 162045 65789
rect 161979 65724 161980 65788
rect 162044 65724 162045 65788
rect 161979 65723 162045 65724
rect 163454 64565 163514 75787
rect 163638 74085 163698 79731
rect 163635 74084 163701 74085
rect 163635 74020 163636 74084
rect 163700 74020 163701 74084
rect 163635 74019 163701 74020
rect 163451 64564 163517 64565
rect 163451 64500 163452 64564
rect 163516 64500 163517 64564
rect 163451 64499 163517 64500
rect 161243 63476 161309 63477
rect 161243 63412 161244 63476
rect 161308 63412 161309 63476
rect 161243 63411 161309 63412
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 78000
rect 164558 72589 164618 79731
rect 166582 79661 166642 81227
rect 174859 81156 174925 81157
rect 174859 81092 174860 81156
rect 174924 81092 174925 81156
rect 174859 81091 174925 81092
rect 166947 81020 167013 81021
rect 166947 80956 166948 81020
rect 167012 80956 167013 81020
rect 166947 80955 167013 80956
rect 166763 79932 166829 79933
rect 166763 79868 166764 79932
rect 166828 79868 166829 79932
rect 166763 79867 166829 79868
rect 166395 79660 166461 79661
rect 166395 79596 166396 79660
rect 166460 79596 166461 79660
rect 166395 79595 166461 79596
rect 166579 79660 166645 79661
rect 166579 79596 166580 79660
rect 166644 79596 166645 79660
rect 166579 79595 166645 79596
rect 164923 78572 164989 78573
rect 164923 78508 164924 78572
rect 164988 78508 164989 78572
rect 164923 78507 164989 78508
rect 164555 72588 164621 72589
rect 164555 72524 164556 72588
rect 164620 72524 164621 72588
rect 164555 72523 164621 72524
rect 164926 65653 164986 78507
rect 165843 78300 165909 78301
rect 165843 78236 165844 78300
rect 165908 78236 165909 78300
rect 165843 78235 165909 78236
rect 165846 70277 165906 78235
rect 166398 75930 166458 79595
rect 166398 75870 166642 75930
rect 165843 70276 165909 70277
rect 165843 70212 165844 70276
rect 165908 70212 165909 70276
rect 165843 70211 165909 70212
rect 166582 67285 166642 75870
rect 166579 67284 166645 67285
rect 166579 67220 166580 67284
rect 166644 67220 166645 67284
rect 166579 67219 166645 67220
rect 164923 65652 164989 65653
rect 164923 65588 164924 65652
rect 164988 65588 164989 65652
rect 164923 65587 164989 65588
rect 166766 63341 166826 79867
rect 166950 79797 167010 80955
rect 169155 80204 169221 80205
rect 169155 80140 169156 80204
rect 169220 80140 169221 80204
rect 169155 80139 169221 80140
rect 167131 79932 167197 79933
rect 167131 79868 167132 79932
rect 167196 79868 167197 79932
rect 167131 79867 167197 79868
rect 167867 79932 167933 79933
rect 167867 79868 167868 79932
rect 167932 79868 167933 79932
rect 167867 79867 167933 79868
rect 168235 79932 168301 79933
rect 168235 79868 168236 79932
rect 168300 79868 168301 79932
rect 168235 79867 168301 79868
rect 166947 79796 167013 79797
rect 166947 79732 166948 79796
rect 167012 79732 167013 79796
rect 166947 79731 167013 79732
rect 167134 78845 167194 79867
rect 167683 79796 167749 79797
rect 167683 79732 167684 79796
rect 167748 79732 167749 79796
rect 167683 79731 167749 79732
rect 167131 78844 167197 78845
rect 167131 78780 167132 78844
rect 167196 78780 167197 78844
rect 167131 78779 167197 78780
rect 167686 71501 167746 79731
rect 167870 78981 167930 79867
rect 168051 79660 168117 79661
rect 168051 79596 168052 79660
rect 168116 79596 168117 79660
rect 168051 79595 168117 79596
rect 167867 78980 167933 78981
rect 167867 78916 167868 78980
rect 167932 78916 167933 78980
rect 167867 78915 167933 78916
rect 167867 78844 167933 78845
rect 167867 78780 167868 78844
rect 167932 78780 167933 78844
rect 167867 78779 167933 78780
rect 167683 71500 167749 71501
rect 167683 71436 167684 71500
rect 167748 71436 167749 71500
rect 167683 71435 167749 71436
rect 167870 67149 167930 78779
rect 167867 67148 167933 67149
rect 167867 67084 167868 67148
rect 167932 67084 167933 67148
rect 167867 67083 167933 67084
rect 166763 63340 166829 63341
rect 166763 63276 166764 63340
rect 166828 63276 166829 63340
rect 166763 63275 166829 63276
rect 168054 63205 168114 79595
rect 168238 78981 168298 79867
rect 168235 78980 168301 78981
rect 168235 78916 168236 78980
rect 168300 78916 168301 78980
rect 168235 78915 168301 78916
rect 168051 63204 168117 63205
rect 168051 63140 168052 63204
rect 168116 63140 168117 63204
rect 168051 63139 168117 63140
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 78000
rect 169158 64701 169218 80139
rect 170075 79932 170141 79933
rect 170075 79868 170076 79932
rect 170140 79868 170141 79932
rect 170075 79867 170141 79868
rect 172283 79932 172349 79933
rect 172283 79868 172284 79932
rect 172348 79868 172349 79932
rect 172283 79867 172349 79868
rect 173019 79932 173085 79933
rect 173019 79868 173020 79932
rect 173084 79868 173085 79932
rect 173019 79867 173085 79868
rect 170078 75989 170138 79867
rect 170627 79796 170693 79797
rect 170627 79732 170628 79796
rect 170692 79732 170693 79796
rect 170627 79731 170693 79732
rect 170811 79796 170877 79797
rect 170811 79732 170812 79796
rect 170876 79732 170877 79796
rect 170811 79731 170877 79732
rect 171547 79796 171613 79797
rect 171547 79732 171548 79796
rect 171612 79732 171613 79796
rect 171547 79731 171613 79732
rect 170630 76530 170690 79731
rect 170814 78981 170874 79731
rect 170811 78980 170877 78981
rect 170811 78916 170812 78980
rect 170876 78916 170877 78980
rect 170811 78915 170877 78916
rect 170811 77892 170877 77893
rect 170811 77828 170812 77892
rect 170876 77828 170877 77892
rect 170811 77827 170877 77828
rect 170814 76941 170874 77827
rect 170811 76940 170877 76941
rect 170811 76876 170812 76940
rect 170876 76876 170877 76940
rect 170811 76875 170877 76876
rect 170630 76470 170874 76530
rect 170627 76124 170693 76125
rect 170627 76060 170628 76124
rect 170692 76060 170693 76124
rect 170627 76059 170693 76060
rect 170075 75988 170141 75989
rect 170075 75924 170076 75988
rect 170140 75924 170141 75988
rect 170075 75923 170141 75924
rect 170630 70005 170690 76059
rect 170814 71790 170874 76470
rect 170814 71730 171058 71790
rect 170627 70004 170693 70005
rect 170627 69940 170628 70004
rect 170692 69940 170693 70004
rect 170627 69939 170693 69940
rect 170998 66877 171058 71730
rect 171550 71365 171610 79731
rect 171731 78572 171797 78573
rect 171731 78508 171732 78572
rect 171796 78508 171797 78572
rect 171731 78507 171797 78508
rect 171734 73949 171794 78507
rect 172286 75989 172346 79867
rect 173022 78165 173082 79867
rect 174862 79797 174922 81091
rect 174859 79796 174925 79797
rect 174859 79732 174860 79796
rect 174924 79732 174925 79796
rect 174859 79731 174925 79732
rect 174675 79388 174741 79389
rect 174675 79324 174676 79388
rect 174740 79324 174741 79388
rect 174675 79323 174741 79324
rect 173019 78164 173085 78165
rect 173019 78100 173020 78164
rect 173084 78100 173085 78164
rect 173019 78099 173085 78100
rect 172283 75988 172349 75989
rect 172283 75924 172284 75988
rect 172348 75924 172349 75988
rect 172283 75923 172349 75924
rect 171731 73948 171797 73949
rect 171731 73884 171732 73948
rect 171796 73884 171797 73948
rect 171731 73883 171797 73884
rect 171547 71364 171613 71365
rect 171547 71300 171548 71364
rect 171612 71300 171613 71364
rect 171547 71299 171613 71300
rect 170995 66876 171061 66877
rect 170995 66812 170996 66876
rect 171060 66812 171061 66876
rect 170995 66811 171061 66812
rect 172794 66454 173414 78000
rect 174678 74357 174738 79323
rect 175046 78029 175106 81771
rect 175227 79932 175293 79933
rect 175227 79868 175228 79932
rect 175292 79868 175293 79932
rect 175227 79867 175293 79868
rect 175043 78028 175109 78029
rect 175043 77964 175044 78028
rect 175108 77964 175109 78028
rect 175043 77963 175109 77964
rect 175230 74550 175290 79867
rect 176702 79525 176762 81907
rect 184795 81700 184861 81701
rect 184795 81636 184796 81700
rect 184860 81636 184861 81700
rect 184795 81635 184861 81636
rect 177251 80612 177317 80613
rect 177251 80548 177252 80612
rect 177316 80548 177317 80612
rect 177251 80547 177317 80548
rect 177254 79797 177314 80547
rect 177251 79796 177317 79797
rect 177251 79732 177252 79796
rect 177316 79732 177317 79796
rect 177251 79731 177317 79732
rect 176699 79524 176765 79525
rect 176699 79460 176700 79524
rect 176764 79460 176765 79524
rect 176699 79459 176765 79460
rect 176515 79388 176581 79389
rect 176515 79324 176516 79388
rect 176580 79324 176581 79388
rect 176515 79323 176581 79324
rect 175046 74490 175290 74550
rect 174675 74356 174741 74357
rect 174675 74292 174676 74356
rect 174740 74292 174741 74356
rect 174675 74291 174741 74292
rect 175046 70141 175106 74490
rect 175043 70140 175109 70141
rect 175043 70076 175044 70140
rect 175108 70076 175109 70140
rect 175043 70075 175109 70076
rect 176518 68509 176578 79323
rect 184798 79253 184858 81635
rect 184795 79252 184861 79253
rect 184795 79188 184796 79252
rect 184860 79188 184861 79252
rect 184795 79187 184861 79188
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176515 68508 176581 68509
rect 176515 68444 176516 68508
rect 176580 68444 176581 68508
rect 176515 68443 176581 68444
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 169155 64700 169221 64701
rect 169155 64636 169156 64700
rect 169220 64636 169221 64700
rect 169155 64635 169221 64636
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 186086 65517 186146 82179
rect 186822 80069 186882 136579
rect 186819 80068 186885 80069
rect 186819 80004 186820 80068
rect 186884 80004 186885 80068
rect 186819 80003 186885 80004
rect 187006 78437 187066 139163
rect 187190 137461 187250 139299
rect 187187 137460 187253 137461
rect 187187 137396 187188 137460
rect 187252 137396 187253 137460
rect 187187 137395 187253 137396
rect 187187 82788 187253 82789
rect 187187 82724 187188 82788
rect 187252 82724 187253 82788
rect 187187 82723 187253 82724
rect 187003 78436 187069 78437
rect 187003 78372 187004 78436
rect 187068 78372 187069 78436
rect 187003 78371 187069 78372
rect 186083 65516 186149 65517
rect 186083 65452 186084 65516
rect 186148 65452 186149 65516
rect 186083 65451 186149 65452
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187190 71773 187250 82723
rect 187187 71772 187253 71773
rect 187187 71708 187188 71772
rect 187252 71708 187253 71772
rect 187187 71707 187253 71708
rect 187374 67557 187434 140115
rect 187555 139772 187621 139773
rect 187555 139708 187556 139772
rect 187620 139708 187621 139772
rect 187555 139707 187621 139708
rect 187558 137325 187618 139707
rect 187555 137324 187621 137325
rect 187555 137260 187556 137324
rect 187620 137260 187621 137324
rect 187555 137259 187621 137260
rect 187742 69869 187802 189619
rect 187923 186964 187989 186965
rect 187923 186900 187924 186964
rect 187988 186900 187989 186964
rect 187923 186899 187989 186900
rect 187739 69868 187805 69869
rect 187739 69804 187740 69868
rect 187804 69804 187805 69868
rect 187739 69803 187805 69804
rect 187926 69461 187986 186899
rect 188107 140044 188173 140045
rect 188107 139980 188108 140044
rect 188172 139980 188173 140044
rect 188107 139979 188173 139980
rect 188110 71093 188170 139979
rect 189030 78029 189090 190707
rect 189211 185604 189277 185605
rect 189211 185540 189212 185604
rect 189276 185540 189277 185604
rect 189211 185539 189277 185540
rect 189214 78165 189274 185539
rect 189211 78164 189277 78165
rect 189211 78100 189212 78164
rect 189276 78100 189277 78164
rect 189211 78099 189277 78100
rect 189027 78028 189093 78029
rect 189027 77964 189028 78028
rect 189092 77964 189093 78028
rect 189027 77963 189093 77964
rect 190502 74221 190562 196555
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 142000 191414 155898
rect 191790 142765 191850 262923
rect 194550 262853 194610 268363
rect 193259 262852 193325 262853
rect 193259 262788 193260 262852
rect 193324 262788 193325 262852
rect 193259 262787 193325 262788
rect 194547 262852 194613 262853
rect 194547 262788 194548 262852
rect 194612 262788 194613 262852
rect 194547 262787 194613 262788
rect 191971 190092 192037 190093
rect 191971 190028 191972 190092
rect 192036 190028 192037 190092
rect 191971 190027 192037 190028
rect 193075 190092 193141 190093
rect 193075 190028 193076 190092
rect 193140 190028 193141 190092
rect 193075 190027 193141 190028
rect 191787 142764 191853 142765
rect 191787 142700 191788 142764
rect 191852 142700 191853 142764
rect 191787 142699 191853 142700
rect 190683 138956 190749 138957
rect 190683 138892 190684 138956
rect 190748 138892 190749 138956
rect 190683 138891 190749 138892
rect 190686 80613 190746 138891
rect 190683 80612 190749 80613
rect 190683 80548 190684 80612
rect 190748 80548 190749 80612
rect 190683 80547 190749 80548
rect 190499 74220 190565 74221
rect 190499 74156 190500 74220
rect 190564 74156 190565 74220
rect 190499 74155 190565 74156
rect 188107 71092 188173 71093
rect 188107 71028 188108 71092
rect 188172 71028 188173 71092
rect 188107 71027 188173 71028
rect 187923 69460 187989 69461
rect 187923 69396 187924 69460
rect 187988 69396 187989 69460
rect 187923 69395 187989 69396
rect 187371 67556 187437 67557
rect 187371 67492 187372 67556
rect 187436 67492 187437 67556
rect 187371 67491 187437 67492
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191974 72453 192034 190027
rect 193078 189685 193138 190027
rect 193075 189684 193141 189685
rect 193075 189620 193076 189684
rect 193140 189620 193141 189684
rect 193075 189619 193141 189620
rect 192155 144124 192221 144125
rect 192155 144060 192156 144124
rect 192220 144060 192221 144124
rect 192155 144059 192221 144060
rect 191971 72452 192037 72453
rect 191971 72388 191972 72452
rect 192036 72388 192037 72452
rect 191971 72387 192037 72388
rect 192158 66741 192218 144059
rect 193262 142901 193322 262787
rect 195294 232954 195914 268398
rect 196022 262581 196082 269723
rect 196203 263668 196269 263669
rect 196203 263604 196204 263668
rect 196268 263604 196269 263668
rect 196203 263603 196269 263604
rect 196019 262580 196085 262581
rect 196019 262516 196020 262580
rect 196084 262516 196085 262580
rect 196019 262515 196085 262516
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 193259 142900 193325 142901
rect 193259 142836 193260 142900
rect 193324 142836 193325 142900
rect 193259 142835 193325 142836
rect 193443 141676 193509 141677
rect 193443 141612 193444 141676
rect 193508 141612 193509 141676
rect 193443 141611 193509 141612
rect 193259 137868 193325 137869
rect 193259 137804 193260 137868
rect 193324 137804 193325 137868
rect 193259 137803 193325 137804
rect 192155 66740 192221 66741
rect 192155 66676 192156 66740
rect 192220 66676 192221 66740
rect 192155 66675 192221 66676
rect 193262 64837 193322 137803
rect 193446 71637 193506 141611
rect 194547 141404 194613 141405
rect 194547 141340 194548 141404
rect 194612 141340 194613 141404
rect 194547 141339 194613 141340
rect 193627 140588 193693 140589
rect 193627 140524 193628 140588
rect 193692 140524 193693 140588
rect 193627 140523 193693 140524
rect 193630 73813 193690 140523
rect 193811 138820 193877 138821
rect 193811 138756 193812 138820
rect 193876 138756 193877 138820
rect 193811 138755 193877 138756
rect 193814 82245 193874 138755
rect 193811 82244 193877 82245
rect 193811 82180 193812 82244
rect 193876 82180 193877 82244
rect 193811 82179 193877 82180
rect 193627 73812 193693 73813
rect 193627 73748 193628 73812
rect 193692 73748 193693 73812
rect 193627 73747 193693 73748
rect 193443 71636 193509 71637
rect 193443 71572 193444 71636
rect 193508 71572 193509 71636
rect 193443 71571 193509 71572
rect 193259 64836 193325 64837
rect 193259 64772 193260 64836
rect 193324 64772 193325 64836
rect 193259 64771 193325 64772
rect 194550 64565 194610 141339
rect 194731 140316 194797 140317
rect 194731 140252 194732 140316
rect 194796 140252 194797 140316
rect 194731 140251 194797 140252
rect 194734 73677 194794 140251
rect 195294 124954 195914 160398
rect 196022 143309 196082 262515
rect 196206 145757 196266 263603
rect 197491 262444 197557 262445
rect 197491 262380 197492 262444
rect 197556 262380 197557 262444
rect 197491 262379 197557 262380
rect 197307 194036 197373 194037
rect 197307 193972 197308 194036
rect 197372 193972 197373 194036
rect 197307 193971 197373 193972
rect 197310 190637 197370 193971
rect 197307 190636 197373 190637
rect 197307 190572 197308 190636
rect 197372 190572 197373 190636
rect 197307 190571 197373 190572
rect 196203 145756 196269 145757
rect 196203 145692 196204 145756
rect 196268 145692 196269 145756
rect 196203 145691 196269 145692
rect 196571 144396 196637 144397
rect 196571 144332 196572 144396
rect 196636 144332 196637 144396
rect 196571 144331 196637 144332
rect 196019 143308 196085 143309
rect 196019 143244 196020 143308
rect 196084 143244 196085 143308
rect 196019 143243 196085 143244
rect 196387 141540 196453 141541
rect 196387 141476 196388 141540
rect 196452 141476 196453 141540
rect 196387 141475 196453 141476
rect 196203 140044 196269 140045
rect 196203 139980 196204 140044
rect 196268 139980 196269 140044
rect 196203 139979 196269 139980
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194731 73676 194797 73677
rect 194731 73612 194732 73676
rect 194796 73612 194797 73676
rect 194731 73611 194797 73612
rect 194547 64564 194613 64565
rect 194547 64500 194548 64564
rect 194612 64500 194613 64564
rect 194547 64499 194613 64500
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 88398
rect 196206 74085 196266 139979
rect 196390 81429 196450 141475
rect 196387 81428 196453 81429
rect 196387 81364 196388 81428
rect 196452 81364 196453 81428
rect 196387 81363 196453 81364
rect 196203 74084 196269 74085
rect 196203 74020 196204 74084
rect 196268 74020 196269 74084
rect 196203 74019 196269 74020
rect 196574 69733 196634 144331
rect 197310 73133 197370 190571
rect 197494 146029 197554 262379
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198779 193900 198845 193901
rect 198779 193836 198780 193900
rect 198844 193836 198845 193900
rect 198779 193835 198845 193836
rect 197491 146028 197557 146029
rect 197491 145964 197492 146028
rect 197556 145964 197557 146028
rect 197491 145963 197557 145964
rect 198782 76669 198842 193835
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200619 192540 200685 192541
rect 200619 192476 200620 192540
rect 200684 192476 200685 192540
rect 200619 192475 200685 192476
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 198963 146980 199029 146981
rect 198963 146916 198964 146980
rect 199028 146916 199029 146980
rect 198963 146915 199029 146916
rect 198779 76668 198845 76669
rect 198779 76604 198780 76668
rect 198844 76604 198845 76668
rect 198779 76603 198845 76604
rect 197307 73132 197373 73133
rect 197307 73068 197308 73132
rect 197372 73068 197373 73132
rect 197307 73067 197373 73068
rect 196571 69732 196637 69733
rect 196571 69668 196572 69732
rect 196636 69668 196637 69732
rect 196571 69667 196637 69668
rect 198966 67421 199026 146915
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198963 67420 199029 67421
rect 198963 67356 198964 67420
rect 199028 67356 199029 67420
rect 198963 67355 199029 67356
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 92898
rect 200622 67013 200682 192475
rect 202091 191588 202157 191589
rect 202091 191524 202092 191588
rect 202156 191524 202157 191588
rect 202091 191523 202157 191524
rect 201539 188460 201605 188461
rect 201539 188396 201540 188460
rect 201604 188396 201605 188460
rect 201539 188395 201605 188396
rect 201542 72861 201602 188395
rect 201539 72860 201605 72861
rect 201539 72796 201540 72860
rect 201604 72796 201605 72860
rect 201539 72795 201605 72796
rect 202094 70277 202154 191523
rect 203563 184244 203629 184245
rect 203563 184180 203564 184244
rect 203628 184180 203629 184244
rect 203563 184179 203629 184180
rect 203011 178804 203077 178805
rect 203011 178740 203012 178804
rect 203076 178740 203077 178804
rect 203011 178739 203077 178740
rect 202091 70276 202157 70277
rect 202091 70212 202092 70276
rect 202156 70212 202157 70276
rect 202091 70211 202157 70212
rect 203014 68645 203074 178739
rect 203566 81157 203626 184179
rect 204294 169954 204914 205398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 207059 201108 207125 201109
rect 207059 201044 207060 201108
rect 207124 201044 207125 201108
rect 207059 201043 207125 201044
rect 205035 200972 205101 200973
rect 205035 200908 205036 200972
rect 205100 200908 205101 200972
rect 205035 200907 205101 200908
rect 205038 200565 205098 200907
rect 205035 200564 205101 200565
rect 205035 200500 205036 200564
rect 205100 200500 205101 200564
rect 205035 200499 205101 200500
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203563 81156 203629 81157
rect 203563 81092 203564 81156
rect 203628 81092 203629 81156
rect 203563 81091 203629 81092
rect 203011 68644 203077 68645
rect 203011 68580 203012 68644
rect 203076 68580 203077 68644
rect 203011 68579 203077 68580
rect 200619 67012 200685 67013
rect 200619 66948 200620 67012
rect 200684 66948 200685 67012
rect 200619 66947 200685 66948
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 61954 204914 97398
rect 205038 70277 205098 200499
rect 207062 200429 207122 201043
rect 207059 200428 207125 200429
rect 207059 200364 207060 200428
rect 207124 200364 207125 200428
rect 207059 200363 207125 200364
rect 205587 199612 205653 199613
rect 205587 199548 205588 199612
rect 205652 199548 205653 199612
rect 205587 199547 205653 199548
rect 205590 198933 205650 199547
rect 205587 198932 205653 198933
rect 205587 198868 205588 198932
rect 205652 198868 205653 198932
rect 205587 198867 205653 198868
rect 206139 198932 206205 198933
rect 206139 198868 206140 198932
rect 206204 198868 206205 198932
rect 206139 198867 206205 198868
rect 205587 196756 205653 196757
rect 205587 196692 205588 196756
rect 205652 196692 205653 196756
rect 205587 196691 205653 196692
rect 205590 71365 205650 196691
rect 205771 193084 205837 193085
rect 205771 193020 205772 193084
rect 205836 193020 205837 193084
rect 205771 193019 205837 193020
rect 205587 71364 205653 71365
rect 205587 71300 205588 71364
rect 205652 71300 205653 71364
rect 205587 71299 205653 71300
rect 205774 71229 205834 193019
rect 205771 71228 205837 71229
rect 205771 71164 205772 71228
rect 205836 71164 205837 71228
rect 205771 71163 205837 71164
rect 205035 70276 205101 70277
rect 205035 70212 205036 70276
rect 205100 70212 205101 70276
rect 205035 70211 205101 70212
rect 206142 70005 206202 198867
rect 207062 70141 207122 200363
rect 207611 187372 207677 187373
rect 207611 187308 207612 187372
rect 207676 187308 207677 187372
rect 207611 187307 207677 187308
rect 207614 71501 207674 187307
rect 208794 174454 209414 209898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 210923 200836 210989 200837
rect 210923 200772 210924 200836
rect 210988 200772 210989 200836
rect 210923 200771 210989 200772
rect 210926 200157 210986 200771
rect 211107 200700 211173 200701
rect 211107 200636 211108 200700
rect 211172 200636 211173 200700
rect 211107 200635 211173 200636
rect 211110 200293 211170 200635
rect 211107 200292 211173 200293
rect 211107 200228 211108 200292
rect 211172 200228 211173 200292
rect 211107 200227 211173 200228
rect 209819 200156 209885 200157
rect 209819 200092 209820 200156
rect 209884 200092 209885 200156
rect 209819 200091 209885 200092
rect 210923 200156 210989 200157
rect 210923 200092 210924 200156
rect 210988 200092 210989 200156
rect 210923 200091 210989 200092
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 207611 71500 207677 71501
rect 207611 71436 207612 71500
rect 207676 71436 207677 71500
rect 207611 71435 207677 71436
rect 207059 70140 207125 70141
rect 207059 70076 207060 70140
rect 207124 70076 207125 70140
rect 207059 70075 207125 70076
rect 206139 70004 206205 70005
rect 206139 69940 206140 70004
rect 206204 69940 206205 70004
rect 206139 69939 206205 69940
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 66454 209414 101898
rect 209822 68509 209882 200091
rect 210371 197028 210437 197029
rect 210371 196964 210372 197028
rect 210436 196964 210437 197028
rect 210371 196963 210437 196964
rect 210923 197028 210989 197029
rect 210923 196964 210924 197028
rect 210988 196964 210989 197028
rect 210923 196963 210989 196964
rect 210374 76805 210434 196963
rect 210926 196757 210986 196963
rect 210923 196756 210989 196757
rect 210923 196692 210924 196756
rect 210988 196692 210989 196756
rect 210923 196691 210989 196692
rect 210371 76804 210437 76805
rect 210371 76740 210372 76804
rect 210436 76740 210437 76804
rect 210371 76739 210437 76740
rect 211110 76669 211170 200227
rect 213294 178954 213914 214398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 214051 195124 214117 195125
rect 214051 195060 214052 195124
rect 214116 195060 214117 195124
rect 214051 195059 214117 195060
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 211107 76668 211173 76669
rect 211107 76604 211108 76668
rect 211172 76604 211173 76668
rect 211107 76603 211173 76604
rect 213294 70954 213914 106398
rect 214054 75445 214114 195059
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 214051 75444 214117 75445
rect 214051 75380 214052 75444
rect 214116 75380 214117 75444
rect 214051 75379 214117 75380
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 209819 68508 209885 68509
rect 209819 68444 209820 68508
rect 209884 68444 209885 68508
rect 209819 68443 209885 68444
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 570 0 69354 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal2 s 87574 -960 87686 480 0 FreeSans 448 90 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal2 s 156482 -960 156594 480 0 FreeSans 448 90 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 583520 56388 584960 56628 0 FreeSans 960 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal2 s 100454 703520 100566 704960 0 FreeSans 448 90 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -960 326348 480 326588 0 FreeSans 960 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal2 s 345174 703520 345286 704960 0 FreeSans 448 90 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s 583520 222308 584960 222548 0 FreeSans 960 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -960 637108 480 637348 0 FreeSans 960 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 128468 480 128708 0 FreeSans 960 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 80868 584960 81108 0 FreeSans 960 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal2 s 259522 -960 259634 480 0 FreeSans 448 90 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s -960 435148 480 435388 0 FreeSans 960 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 673828 584960 674068 0 FreeSans 960 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s -960 205308 480 205548 0 FreeSans 960 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s -960 399108 480 399348 0 FreeSans 960 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal2 s 75982 -960 76094 480 0 FreeSans 448 90 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal2 s 546102 -960 546214 480 0 FreeSans 448 90 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal2 s 412150 -960 412262 480 0 FreeSans 448 90 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal2 s 240202 -960 240314 480 0 FreeSans 448 90 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -960 536468 480 536708 0 FreeSans 960 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -960 447388 480 447628 0 FreeSans 960 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal2 s 173226 703520 173338 704960 0 FreeSans 448 90 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal2 s 390898 703520 391010 704960 0 FreeSans 448 90 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -960 382788 480 383028 0 FreeSans 960 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -960 59788 480 60028 0 FreeSans 960 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s 583520 28508 584960 28748 0 FreeSans 960 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal2 s 211222 703520 211334 704960 0 FreeSans 448 90 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal2 s 121706 -960 121818 480 0 FreeSans 448 90 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal2 s 328430 -960 328542 480 0 FreeSans 448 90 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 641868 584960 642108 0 FreeSans 960 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal2 s 191902 703520 192014 704960 0 FreeSans 448 90 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 64548 584960 64788 0 FreeSans 960 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 601068 584960 601308 0 FreeSans 960 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 583520 492268 584960 492508 0 FreeSans 960 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -960 88348 480 88588 0 FreeSans 960 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -960 132548 480 132788 0 FreeSans 960 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s -960 245428 480 245668 0 FreeSans 960 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal2 s 56662 -960 56774 480 0 FreeSans 448 90 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 583520 60468 584960 60708 0 FreeSans 960 0 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 583520 552788 584960 553028 0 FreeSans 960 0 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal2 s 228610 -960 228722 480 0 FreeSans 448 90 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal2 s 88862 703520 88974 704960 0 FreeSans 448 90 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal2 s 450790 -960 450902 480 0 FreeSans 448 90 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s -960 233868 480 234108 0 FreeSans 960 0 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal2 s 209934 -960 210046 480 0 FreeSans 448 90 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s -960 334508 480 334748 0 FreeSans 960 0 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal2 s 22530 -960 22642 480 0 FreeSans 448 90 0 0 io_clamp_high[0]
port 47 nsew signal bidirectional
flabel metal3 s 583520 581348 584960 581588 0 FreeSans 960 0 0 0 io_clamp_high[1]
port 48 nsew signal bidirectional
flabel metal3 s 583520 363068 584960 363308 0 FreeSans 960 0 0 0 io_clamp_high[2]
port 49 nsew signal bidirectional
flabel metal3 s -960 124388 480 124628 0 FreeSans 960 0 0 0 io_clamp_low[0]
port 50 nsew signal bidirectional
flabel metal2 s 285926 -960 286038 480 0 FreeSans 448 90 0 0 io_clamp_low[1]
port 51 nsew signal bidirectional
flabel metal3 s -960 649348 480 649588 0 FreeSans 960 0 0 0 io_clamp_low[2]
port 52 nsew signal bidirectional
flabel metal2 s 37986 -960 38098 480 0 FreeSans 448 90 0 0 io_in[0]
port 53 nsew signal input
flabel metal3 s 583520 504508 584960 504748 0 FreeSans 960 0 0 0 io_in[10]
port 54 nsew signal input
flabel metal2 s 493938 703520 494050 704960 0 FreeSans 448 90 0 0 io_in[11]
port 55 nsew signal input
flabel metal2 s 402490 703520 402602 704960 0 FreeSans 448 90 0 0 io_in[12]
port 56 nsew signal input
flabel metal2 s 99166 -960 99278 480 0 FreeSans 448 90 0 0 io_in[13]
port 57 nsew signal input
flabel metal2 s 416014 -960 416126 480 0 FreeSans 448 90 0 0 io_in[14]
port 58 nsew signal input
flabel metal3 s -960 76108 480 76348 0 FreeSans 960 0 0 0 io_in[15]
port 59 nsew signal input
flabel metal2 s 519054 -960 519166 480 0 FreeSans 448 90 0 0 io_in[16]
port 60 nsew signal input
flabel metal3 s 583520 237948 584960 238188 0 FreeSans 960 0 0 0 io_in[17]
port 61 nsew signal input
flabel metal3 s 583520 72708 584960 72948 0 FreeSans 960 0 0 0 io_in[18]
port 62 nsew signal input
flabel metal3 s -960 564348 480 564588 0 FreeSans 960 0 0 0 io_in[19]
port 63 nsew signal input
flabel metal2 s 492650 -960 492762 480 0 FreeSans 448 90 0 0 io_in[1]
port 64 nsew signal input
flabel metal2 s 534510 -960 534622 480 0 FreeSans 448 90 0 0 io_in[20]
port 65 nsew signal input
flabel metal2 s 336158 -960 336270 480 0 FreeSans 448 90 0 0 io_in[21]
port 66 nsew signal input
flabel metal3 s 583520 133228 584960 133468 0 FreeSans 960 0 0 0 io_in[22]
port 67 nsew signal input
flabel metal2 s 264674 703520 264786 704960 0 FreeSans 448 90 0 0 io_in[23]
port 68 nsew signal input
flabel metal3 s 583520 399788 584960 400028 0 FreeSans 960 0 0 0 io_in[24]
port 69 nsew signal input
flabel metal2 s 580234 -960 580346 480 0 FreeSans 448 90 0 0 io_in[25]
port 70 nsew signal input
flabel metal2 s 535798 703520 535910 704960 0 FreeSans 448 90 0 0 io_in[26]
port 71 nsew signal input
flabel metal3 s 583520 452148 584960 452388 0 FreeSans 960 0 0 0 io_in[2]
port 72 nsew signal input
flabel metal3 s -960 314108 480 314348 0 FreeSans 960 0 0 0 io_in[3]
port 73 nsew signal input
flabel metal2 s 427606 -960 427718 480 0 FreeSans 448 90 0 0 io_in[4]
port 74 nsew signal input
flabel metal2 s 130722 703520 130834 704960 0 FreeSans 448 90 0 0 io_in[5]
port 75 nsew signal input
flabel metal3 s 583520 548708 584960 548948 0 FreeSans 960 0 0 0 io_in[6]
port 76 nsew signal input
flabel metal3 s -960 56388 480 56628 0 FreeSans 960 0 0 0 io_in[7]
port 77 nsew signal input
flabel metal2 s 83710 -960 83822 480 0 FreeSans 448 90 0 0 io_in[8]
port 78 nsew signal input
flabel metal2 s 230542 703520 230654 704960 0 FreeSans 448 90 0 0 io_in[9]
port 79 nsew signal input
flabel metal2 s 164210 -960 164322 480 0 FreeSans 448 90 0 0 io_in_3v3[0]
port 80 nsew signal input
flabel metal2 s 45714 -960 45826 480 0 FreeSans 448 90 0 0 io_in_3v3[10]
port 81 nsew signal input
flabel metal2 s 337446 703520 337558 704960 0 FreeSans 448 90 0 0 io_in_3v3[11]
port 82 nsew signal input
flabel metal2 s 531934 703520 532046 704960 0 FreeSans 448 90 0 0 io_in_3v3[12]
port 83 nsew signal input
flabel metal2 s 10938 -960 11050 480 0 FreeSans 448 90 0 0 io_in_3v3[13]
port 84 nsew signal input
flabel metal3 s -960 641188 480 641428 0 FreeSans 960 0 0 0 io_in_3v3[14]
port 85 nsew signal input
flabel metal3 s 583520 205988 584960 206228 0 FreeSans 960 0 0 0 io_in_3v3[15]
port 86 nsew signal input
flabel metal3 s 583520 157708 584960 157948 0 FreeSans 960 0 0 0 io_in_3v3[16]
port 87 nsew signal input
flabel metal3 s -960 657508 480 657748 0 FreeSans 960 0 0 0 io_in_3v3[17]
port 88 nsew signal input
flabel metal3 s -960 366468 480 366708 0 FreeSans 960 0 0 0 io_in_3v3[18]
port 89 nsew signal input
flabel metal3 s -960 633028 480 633268 0 FreeSans 960 0 0 0 io_in_3v3[19]
port 90 nsew signal input
flabel metal3 s 583520 52308 584960 52548 0 FreeSans 960 0 0 0 io_in_3v3[1]
port 91 nsew signal input
flabel metal2 s 73406 703520 73518 704960 0 FreeSans 448 90 0 0 io_in_3v3[20]
port 92 nsew signal input
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 io_in_3v3[21]
port 93 nsew signal input
flabel metal3 s -960 697628 480 697868 0 FreeSans 960 0 0 0 io_in_3v3[22]
port 94 nsew signal input
flabel metal3 s -960 677228 480 677468 0 FreeSans 960 0 0 0 io_in_3v3[23]
port 95 nsew signal input
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 io_in_3v3[24]
port 96 nsew signal input
flabel metal3 s 583520 335188 584960 335428 0 FreeSans 960 0 0 0 io_in_3v3[25]
port 97 nsew signal input
flabel metal3 s -960 395028 480 395268 0 FreeSans 960 0 0 0 io_in_3v3[26]
port 98 nsew signal input
flabel metal2 s 1278 703520 1390 704960 0 FreeSans 448 90 0 0 io_in_3v3[2]
port 99 nsew signal input
flabel metal3 s 583520 653428 584960 653668 0 FreeSans 960 0 0 0 io_in_3v3[3]
port 100 nsew signal input
flabel metal2 s 566710 703520 566822 704960 0 FreeSans 448 90 0 0 io_in_3v3[4]
port 101 nsew signal input
flabel metal2 s 312974 -960 313086 480 0 FreeSans 448 90 0 0 io_in_3v3[5]
port 102 nsew signal input
flabel metal2 s 446926 -960 447038 480 0 FreeSans 448 90 0 0 io_in_3v3[6]
port 103 nsew signal input
flabel metal2 s 198342 -960 198454 480 0 FreeSans 448 90 0 0 io_in_3v3[7]
port 104 nsew signal input
flabel metal2 s 295586 703520 295698 704960 0 FreeSans 448 90 0 0 io_in_3v3[8]
port 105 nsew signal input
flabel metal2 s 553830 -960 553942 480 0 FreeSans 448 90 0 0 io_in_3v3[9]
port 106 nsew signal input
flabel metal3 s -960 475948 480 476188 0 FreeSans 960 0 0 0 io_oeb[0]
port 107 nsew signal tristate
flabel metal2 s 474618 703520 474730 704960 0 FreeSans 448 90 0 0 io_oeb[10]
port 108 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_oeb[11]
port 109 nsew signal tristate
flabel metal2 s 366426 -960 366538 480 0 FreeSans 448 90 0 0 io_oeb[12]
port 110 nsew signal tristate
flabel metal2 s 515190 -960 515302 480 0 FreeSans 448 90 0 0 io_oeb[13]
port 111 nsew signal tristate
flabel metal3 s 583520 350828 584960 351068 0 FreeSans 960 0 0 0 io_oeb[14]
port 112 nsew signal tristate
flabel metal3 s -960 487508 480 487748 0 FreeSans 960 0 0 0 io_oeb[15]
port 113 nsew signal tristate
flabel metal3 s -960 528308 480 528548 0 FreeSans 960 0 0 0 io_oeb[16]
port 114 nsew signal tristate
flabel metal3 s 583520 592908 584960 593148 0 FreeSans 960 0 0 0 io_oeb[17]
port 115 nsew signal tristate
flabel metal2 s 129434 -960 129546 480 0 FreeSans 448 90 0 0 io_oeb[18]
port 116 nsew signal tristate
flabel metal3 s 583520 649348 584960 649588 0 FreeSans 960 0 0 0 io_oeb[19]
port 117 nsew signal tristate
flabel metal2 s 501666 703520 501778 704960 0 FreeSans 448 90 0 0 io_oeb[1]
port 118 nsew signal tristate
flabel metal2 s 524850 703520 524962 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 119 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 120 nsew signal tristate
flabel metal2 s 60526 -960 60638 480 0 FreeSans 448 90 0 0 io_oeb[22]
port 121 nsew signal tristate
flabel metal3 s 583520 169268 584960 169508 0 FreeSans 960 0 0 0 io_oeb[23]
port 122 nsew signal tristate
flabel metal2 s 349038 703520 349150 704960 0 FreeSans 448 90 0 0 io_oeb[24]
port 123 nsew signal tristate
flabel metal3 s 583520 484108 584960 484348 0 FreeSans 960 0 0 0 io_oeb[25]
port 124 nsew signal tristate
flabel metal3 s 583520 375308 584960 375548 0 FreeSans 960 0 0 0 io_oeb[26]
port 125 nsew signal tristate
flabel metal3 s -960 608548 480 608788 0 FreeSans 960 0 0 0 io_oeb[2]
port 126 nsew signal tristate
flabel metal3 s -960 624868 480 625108 0 FreeSans 960 0 0 0 io_oeb[3]
port 127 nsew signal tristate
flabel metal3 s -960 467788 480 468028 0 FreeSans 960 0 0 0 io_oeb[4]
port 128 nsew signal tristate
flabel metal3 s 583520 560948 584960 561188 0 FreeSans 960 0 0 0 io_oeb[5]
port 129 nsew signal tristate
flabel metal2 s 39274 703520 39386 704960 0 FreeSans 448 90 0 0 io_oeb[6]
port 130 nsew signal tristate
flabel metal3 s -960 520148 480 520388 0 FreeSans 960 0 0 0 io_oeb[7]
port 131 nsew signal tristate
flabel metal2 s 299450 703520 299562 704960 0 FreeSans 448 90 0 0 io_oeb[8]
port 132 nsew signal tristate
flabel metal3 s 583520 294388 584960 294628 0 FreeSans 960 0 0 0 io_oeb[9]
port 133 nsew signal tristate
flabel metal2 s 520986 703520 521098 704960 0 FreeSans 448 90 0 0 io_out[0]
port 134 nsew signal tristate
flabel metal3 s -960 177428 480 177668 0 FreeSans 960 0 0 0 io_out[10]
port 135 nsew signal tristate
flabel metal3 s 583520 665668 584960 665908 0 FreeSans 960 0 0 0 io_out[11]
port 136 nsew signal tristate
flabel metal3 s -960 298468 480 298708 0 FreeSans 960 0 0 0 io_out[12]
port 137 nsew signal tristate
flabel metal3 s 583520 415428 584960 415668 0 FreeSans 960 0 0 0 io_out[13]
port 138 nsew signal tristate
flabel metal2 s 268538 703520 268650 704960 0 FreeSans 448 90 0 0 io_out[14]
port 139 nsew signal tristate
flabel metal3 s -960 346748 480 346988 0 FreeSans 960 0 0 0 io_out[15]
port 140 nsew signal tristate
flabel metal2 s 58594 703520 58706 704960 0 FreeSans 448 90 0 0 io_out[16]
port 141 nsew signal tristate
flabel metal2 s 195766 703520 195878 704960 0 FreeSans 448 90 0 0 io_out[17]
port 142 nsew signal tristate
flabel metal2 s 23818 703520 23930 704960 0 FreeSans 448 90 0 0 io_out[18]
port 143 nsew signal tristate
flabel metal3 s 583520 266508 584960 266748 0 FreeSans 960 0 0 0 io_out[19]
port 144 nsew signal tristate
flabel metal3 s 583520 407268 584960 407508 0 FreeSans 960 0 0 0 io_out[1]
port 145 nsew signal tristate
flabel metal2 s 70186 703520 70298 704960 0 FreeSans 448 90 0 0 io_out[20]
port 146 nsew signal tristate
flabel metal2 s 271114 -960 271226 480 0 FreeSans 448 90 0 0 io_out[21]
port 147 nsew signal tristate
flabel metal3 s -960 184908 480 185148 0 FreeSans 960 0 0 0 io_out[22]
port 148 nsew signal tristate
flabel metal3 s 583520 354908 584960 355148 0 FreeSans 960 0 0 0 io_out[23]
port 149 nsew signal tristate
flabel metal3 s -960 685388 480 685628 0 FreeSans 960 0 0 0 io_out[24]
port 150 nsew signal tristate
flabel metal3 s -960 269908 480 270148 0 FreeSans 960 0 0 0 io_out[25]
port 151 nsew signal tristate
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 io_out[26]
port 152 nsew signal tristate
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 io_out[2]
port 153 nsew signal tristate
flabel metal2 s 276266 703520 276378 704960 0 FreeSans 448 90 0 0 io_out[3]
port 154 nsew signal tristate
flabel metal2 s 470754 703520 470866 704960 0 FreeSans 448 90 0 0 io_out[4]
port 155 nsew signal tristate
flabel metal3 s -960 483428 480 483668 0 FreeSans 960 0 0 0 io_out[5]
port 156 nsew signal tristate
flabel metal3 s 583520 165188 584960 165428 0 FreeSans 960 0 0 0 io_out[6]
port 157 nsew signal tristate
flabel metal3 s -960 653428 480 653668 0 FreeSans 960 0 0 0 io_out[7]
port 158 nsew signal tristate
flabel metal3 s 583520 120988 584960 121228 0 FreeSans 960 0 0 0 io_out[8]
port 159 nsew signal tristate
flabel metal3 s 583520 250188 584960 250428 0 FreeSans 960 0 0 0 io_out[9]
port 160 nsew signal tristate
flabel metal2 s 157770 703520 157882 704960 0 FreeSans 448 90 0 0 la_data_in[0]
port 161 nsew signal input
flabel metal3 s 583520 625548 584960 625788 0 FreeSans 960 0 0 0 la_data_in[100]
port 162 nsew signal input
flabel metal3 s 583520 214148 584960 214388 0 FreeSans 960 0 0 0 la_data_in[101]
port 163 nsew signal input
flabel metal2 s 387034 703520 387146 704960 0 FreeSans 448 90 0 0 la_data_in[102]
port 164 nsew signal input
flabel metal3 s 583520 20348 584960 20588 0 FreeSans 960 0 0 0 la_data_in[103]
port 165 nsew signal input
flabel metal3 s -960 370548 480 370788 0 FreeSans 960 0 0 0 la_data_in[104]
port 166 nsew signal input
flabel metal2 s 222814 703520 222926 704960 0 FreeSans 448 90 0 0 la_data_in[105]
port 167 nsew signal input
flabel metal2 s 134586 703520 134698 704960 0 FreeSans 448 90 0 0 la_data_in[106]
port 168 nsew signal input
flabel metal3 s -960 415428 480 415668 0 FreeSans 960 0 0 0 la_data_in[107]
port 169 nsew signal input
flabel metal3 s 583520 584748 584960 584988 0 FreeSans 960 0 0 0 la_data_in[108]
port 170 nsew signal input
flabel metal3 s -960 161108 480 161348 0 FreeSans 960 0 0 0 la_data_in[109]
port 171 nsew signal input
flabel metal3 s 583520 379388 584960 379628 0 FreeSans 960 0 0 0 la_data_in[10]
port 172 nsew signal input
flabel metal3 s -960 286228 480 286468 0 FreeSans 960 0 0 0 la_data_in[110]
port 173 nsew signal input
flabel metal3 s 583520 270588 584960 270828 0 FreeSans 960 0 0 0 la_data_in[111]
port 174 nsew signal input
flabel metal3 s -960 374628 480 374868 0 FreeSans 960 0 0 0 la_data_in[112]
port 175 nsew signal input
flabel metal3 s -960 673148 480 673388 0 FreeSans 960 0 0 0 la_data_in[113]
port 176 nsew signal input
flabel metal3 s -960 516068 480 516308 0 FreeSans 960 0 0 0 la_data_in[114]
port 177 nsew signal input
flabel metal2 s 325854 703520 325966 704960 0 FreeSans 448 90 0 0 la_data_in[115]
port 178 nsew signal input
flabel metal2 s 526782 -960 526894 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 179 nsew signal input
flabel metal3 s -960 338588 480 338828 0 FreeSans 960 0 0 0 la_data_in[117]
port 180 nsew signal input
flabel metal3 s 583520 520828 584960 521068 0 FreeSans 960 0 0 0 la_data_in[118]
port 181 nsew signal input
flabel metal3 s 583520 210068 584960 210308 0 FreeSans 960 0 0 0 la_data_in[119]
port 182 nsew signal input
flabel metal2 s 96590 703520 96702 704960 0 FreeSans 448 90 0 0 la_data_in[11]
port 183 nsew signal input
flabel metal3 s -960 305948 480 306188 0 FreeSans 960 0 0 0 la_data_in[120]
port 184 nsew signal input
flabel metal2 s 160346 -960 160458 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 185 nsew signal input
flabel metal2 s 137162 -960 137274 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 186 nsew signal input
flabel metal3 s -960 426988 480 427228 0 FreeSans 960 0 0 0 la_data_in[123]
port 187 nsew signal input
flabel metal2 s 413438 703520 413550 704960 0 FreeSans 448 90 0 0 la_data_in[124]
port 188 nsew signal input
flabel metal2 s 484922 -960 485034 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 189 nsew signal input
flabel metal3 s -960 419508 480 419748 0 FreeSans 960 0 0 0 la_data_in[126]
port 190 nsew signal input
flabel metal2 s 558982 703520 559094 704960 0 FreeSans 448 90 0 0 la_data_in[127]
port 191 nsew signal input
flabel metal3 s 583520 185588 584960 185828 0 FreeSans 960 0 0 0 la_data_in[12]
port 192 nsew signal input
flabel metal3 s 583520 339268 584960 339508 0 FreeSans 960 0 0 0 la_data_in[13]
port 193 nsew signal input
flabel metal3 s -960 539868 480 540108 0 FreeSans 960 0 0 0 la_data_in[14]
port 194 nsew signal input
flabel metal3 s -960 548028 480 548268 0 FreeSans 960 0 0 0 la_data_in[15]
port 195 nsew signal input
flabel metal3 s -960 67948 480 68188 0 FreeSans 960 0 0 0 la_data_in[16]
port 196 nsew signal input
flabel metal3 s -960 157028 480 157268 0 FreeSans 960 0 0 0 la_data_in[17]
port 197 nsew signal input
flabel metal3 s -960 451468 480 451708 0 FreeSans 960 0 0 0 la_data_in[18]
port 198 nsew signal input
flabel metal2 s 448214 703520 448326 704960 0 FreeSans 448 90 0 0 la_data_in[19]
port 199 nsew signal input
flabel metal2 s 301382 -960 301494 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 200 nsew signal input
flabel metal3 s -960 310028 480 310268 0 FreeSans 960 0 0 0 la_data_in[20]
port 201 nsew signal input
flabel metal2 s 27682 703520 27794 704960 0 FreeSans 448 90 0 0 la_data_in[21]
port 202 nsew signal input
flabel metal2 s 180954 703520 181066 704960 0 FreeSans 448 90 0 0 la_data_in[22]
port 203 nsew signal input
flabel metal3 s -960 439228 480 439468 0 FreeSans 960 0 0 0 la_data_in[23]
port 204 nsew signal input
flabel metal3 s 583520 423588 584960 423828 0 FreeSans 960 0 0 0 la_data_in[24]
port 205 nsew signal input
flabel metal2 s 432758 703520 432870 704960 0 FreeSans 448 90 0 0 la_data_in[25]
port 206 nsew signal input
flabel metal2 s 504242 -960 504354 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 207 nsew signal input
flabel metal2 s 289790 -960 289902 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 208 nsew signal input
flabel metal3 s -960 463708 480 463948 0 FreeSans 960 0 0 0 la_data_in[28]
port 209 nsew signal input
flabel metal3 s -960 342668 480 342908 0 FreeSans 960 0 0 0 la_data_in[29]
port 210 nsew signal input
flabel metal2 s 439198 -960 439310 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 211 nsew signal input
flabel metal3 s -960 491588 480 491828 0 FreeSans 960 0 0 0 la_data_in[30]
port 212 nsew signal input
flabel metal3 s 583520 605148 584960 605388 0 FreeSans 960 0 0 0 la_data_in[31]
port 213 nsew signal input
flabel metal2 s 302670 703520 302782 704960 0 FreeSans 448 90 0 0 la_data_in[32]
port 214 nsew signal input
flabel metal3 s 583520 588828 584960 589068 0 FreeSans 960 0 0 0 la_data_in[33]
port 215 nsew signal input
flabel metal3 s -960 7428 480 7668 0 FreeSans 960 0 0 0 la_data_in[34]
port 216 nsew signal input
flabel metal3 s -960 664988 480 665228 0 FreeSans 960 0 0 0 la_data_in[35]
port 217 nsew signal input
flabel metal2 s 551254 703520 551366 704960 0 FreeSans 448 90 0 0 la_data_in[36]
port 218 nsew signal input
flabel metal2 s 543526 703520 543638 704960 0 FreeSans 448 90 0 0 la_data_in[37]
port 219 nsew signal input
flabel metal2 s 329718 703520 329830 704960 0 FreeSans 448 90 0 0 la_data_in[38]
port 220 nsew signal input
flabel metal2 s 148754 -960 148866 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 221 nsew signal input
flabel metal3 s 583520 395708 584960 395948 0 FreeSans 960 0 0 0 la_data_in[3]
port 222 nsew signal input
flabel metal2 s 138450 703520 138562 704960 0 FreeSans 448 90 0 0 la_data_in[40]
port 223 nsew signal input
flabel metal3 s -960 620788 480 621028 0 FreeSans 960 0 0 0 la_data_in[41]
port 224 nsew signal input
flabel metal3 s -960 144788 480 145028 0 FreeSans 960 0 0 0 la_data_in[42]
port 225 nsew signal input
flabel metal3 s 583520 318868 584960 319108 0 FreeSans 960 0 0 0 la_data_in[43]
port 226 nsew signal input
flabel metal3 s -960 459628 480 459868 0 FreeSans 960 0 0 0 la_data_in[44]
port 227 nsew signal input
flabel metal2 s 81134 703520 81246 704960 0 FreeSans 448 90 0 0 la_data_in[45]
port 228 nsew signal input
flabel metal2 s 123638 703520 123750 704960 0 FreeSans 448 90 0 0 la_data_in[46]
port 229 nsew signal input
flabel metal3 s -960 580668 480 580908 0 FreeSans 960 0 0 0 la_data_in[47]
port 230 nsew signal input
flabel metal3 s 583520 419508 584960 419748 0 FreeSans 960 0 0 0 la_data_in[48]
port 231 nsew signal input
flabel metal3 s 583520 32588 584960 32828 0 FreeSans 960 0 0 0 la_data_in[49]
port 232 nsew signal input
flabel metal2 s 431470 -960 431582 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 233 nsew signal input
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 234 nsew signal input
flabel metal3 s 583520 500428 584960 500668 0 FreeSans 960 0 0 0 la_data_in[51]
port 235 nsew signal input
flabel metal3 s -960 552108 480 552348 0 FreeSans 960 0 0 0 la_data_in[52]
port 236 nsew signal input
flabel metal2 s 255658 -960 255770 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 237 nsew signal input
flabel metal2 s 3210 -960 3322 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 238 nsew signal input
flabel metal3 s 583520 322948 584960 323188 0 FreeSans 960 0 0 0 la_data_in[55]
port 239 nsew signal input
flabel metal3 s -960 507908 480 508148 0 FreeSans 960 0 0 0 la_data_in[56]
port 240 nsew signal input
flabel metal3 s 583520 411348 584960 411588 0 FreeSans 960 0 0 0 la_data_in[57]
port 241 nsew signal input
flabel metal2 s 394762 703520 394874 704960 0 FreeSans 448 90 0 0 la_data_in[58]
port 242 nsew signal input
flabel metal3 s -960 104668 480 104908 0 FreeSans 960 0 0 0 la_data_in[59]
port 243 nsew signal input
flabel metal3 s -960 612628 480 612868 0 FreeSans 960 0 0 0 la_data_in[5]
port 244 nsew signal input
flabel metal2 s 542238 -960 542350 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 245 nsew signal input
flabel metal2 s 568642 -960 568754 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 246 nsew signal input
flabel metal3 s 583520 48228 584960 48468 0 FreeSans 960 0 0 0 la_data_in[62]
port 247 nsew signal input
flabel metal3 s -960 188988 480 189228 0 FreeSans 960 0 0 0 la_data_in[63]
port 248 nsew signal input
flabel metal3 s 583520 173348 584960 173588 0 FreeSans 960 0 0 0 la_data_in[64]
port 249 nsew signal input
flabel metal3 s 583520 577268 584960 577508 0 FreeSans 960 0 0 0 la_data_in[65]
port 250 nsew signal input
flabel metal3 s 583520 331108 584960 331348 0 FreeSans 960 0 0 0 la_data_in[66]
port 251 nsew signal input
flabel metal2 s 79846 -960 79958 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 252 nsew signal input
flabel metal3 s 583520 565028 584960 565268 0 FreeSans 960 0 0 0 la_data_in[68]
port 253 nsew signal input
flabel metal3 s 583520 677908 584960 678148 0 FreeSans 960 0 0 0 la_data_in[69]
port 254 nsew signal input
flabel metal3 s 583520 298468 584960 298708 0 FreeSans 960 0 0 0 la_data_in[6]
port 255 nsew signal input
flabel metal3 s -960 499748 480 499988 0 FreeSans 960 0 0 0 la_data_in[70]
port 256 nsew signal input
flabel metal3 s -960 165188 480 165428 0 FreeSans 960 0 0 0 la_data_in[71]
port 257 nsew signal input
flabel metal2 s 62458 703520 62570 704960 0 FreeSans 448 90 0 0 la_data_in[72]
port 258 nsew signal input
flabel metal3 s -960 100588 480 100828 0 FreeSans 960 0 0 0 la_data_in[73]
port 259 nsew signal input
flabel metal3 s 583520 327028 584960 327268 0 FreeSans 960 0 0 0 la_data_in[74]
port 260 nsew signal input
flabel metal2 s 127502 703520 127614 704960 0 FreeSans 448 90 0 0 la_data_in[75]
port 261 nsew signal input
flabel metal3 s 583520 149548 584960 149788 0 FreeSans 960 0 0 0 la_data_in[76]
port 262 nsew signal input
flabel metal2 s 165498 703520 165610 704960 0 FreeSans 448 90 0 0 la_data_in[77]
port 263 nsew signal input
flabel metal2 s 238270 703520 238382 704960 0 FreeSans 448 90 0 0 la_data_in[78]
port 264 nsew signal input
flabel metal3 s 583520 536468 584960 536708 0 FreeSans 960 0 0 0 la_data_in[79]
port 265 nsew signal input
flabel metal2 s 343242 -960 343354 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 266 nsew signal input
flabel metal3 s -960 330428 480 330668 0 FreeSans 960 0 0 0 la_data_in[80]
port 267 nsew signal input
flabel metal2 s 505530 703520 505642 704960 0 FreeSans 448 90 0 0 la_data_in[81]
port 268 nsew signal input
flabel metal2 s 150042 703520 150154 704960 0 FreeSans 448 90 0 0 la_data_in[82]
port 269 nsew signal input
flabel metal3 s 583520 661588 584960 661828 0 FreeSans 960 0 0 0 la_data_in[83]
port 270 nsew signal input
flabel metal3 s -960 681308 480 681548 0 FreeSans 960 0 0 0 la_data_in[84]
port 271 nsew signal input
flabel metal3 s 583520 367148 584960 367388 0 FreeSans 960 0 0 0 la_data_in[85]
port 272 nsew signal input
flabel metal3 s 583520 448068 584960 448308 0 FreeSans 960 0 0 0 la_data_in[86]
port 273 nsew signal input
flabel metal2 s 95302 -960 95414 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 274 nsew signal input
flabel metal3 s 583520 488188 584960 488428 0 FreeSans 960 0 0 0 la_data_in[88]
port 275 nsew signal input
flabel metal2 s 251794 -960 251906 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 276 nsew signal input
flabel metal2 s 274978 -960 275090 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 277 nsew signal input
flabel metal3 s -960 604468 480 604708 0 FreeSans 960 0 0 0 la_data_in[90]
port 278 nsew signal input
flabel metal3 s -960 532388 480 532628 0 FreeSans 960 0 0 0 la_data_in[91]
port 279 nsew signal input
flabel metal3 s 583520 12188 584960 12428 0 FreeSans 960 0 0 0 la_data_in[92]
port 280 nsew signal input
flabel metal3 s -960 197148 480 197388 0 FreeSans 960 0 0 0 la_data_in[93]
port 281 nsew signal input
flabel metal3 s 583520 314788 584960 315028 0 FreeSans 960 0 0 0 la_data_in[94]
port 282 nsew signal input
flabel metal3 s -960 96508 480 96748 0 FreeSans 960 0 0 0 la_data_in[95]
port 283 nsew signal input
flabel metal3 s -960 511988 480 512228 0 FreeSans 960 0 0 0 la_data_in[96]
port 284 nsew signal input
flabel metal3 s -960 568428 480 568668 0 FreeSans 960 0 0 0 la_data_in[97]
port 285 nsew signal input
flabel metal2 s 282706 -960 282818 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 286 nsew signal input
flabel metal3 s 583520 573188 584960 573428 0 FreeSans 960 0 0 0 la_data_in[99]
port 287 nsew signal input
flabel metal2 s 119774 703520 119886 704960 0 FreeSans 448 90 0 0 la_data_in[9]
port 288 nsew signal input
flabel metal3 s -960 503828 480 504068 0 FreeSans 960 0 0 0 la_data_out[0]
port 289 nsew signal tristate
flabel metal2 s 253082 703520 253194 704960 0 FreeSans 448 90 0 0 la_data_out[100]
port 290 nsew signal tristate
flabel metal2 s 232474 -960 232586 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 291 nsew signal tristate
flabel metal2 s 169362 703520 169474 704960 0 FreeSans 448 90 0 0 la_data_out[102]
port 292 nsew signal tristate
flabel metal3 s 583520 254268 584960 254508 0 FreeSans 960 0 0 0 la_data_out[103]
port 293 nsew signal tristate
flabel metal2 s 161634 703520 161746 704960 0 FreeSans 448 90 0 0 la_data_out[104]
port 294 nsew signal tristate
flabel metal3 s 583520 189668 584960 189908 0 FreeSans 960 0 0 0 la_data_out[105]
port 295 nsew signal tristate
flabel metal2 s 152618 -960 152730 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 296 nsew signal tristate
flabel metal3 s 583520 387548 584960 387788 0 FreeSans 960 0 0 0 la_data_out[107]
port 297 nsew signal tristate
flabel metal3 s 583520 512668 584960 512908 0 FreeSans 960 0 0 0 la_data_out[108]
port 298 nsew signal tristate
flabel metal2 s 509394 703520 509506 704960 0 FreeSans 448 90 0 0 la_data_out[109]
port 299 nsew signal tristate
flabel metal3 s -960 386868 480 387108 0 FreeSans 960 0 0 0 la_data_out[10]
port 300 nsew signal tristate
flabel metal3 s -960 213468 480 213708 0 FreeSans 960 0 0 0 la_data_out[110]
port 301 nsew signal tristate
flabel metal3 s -960 282148 480 282388 0 FreeSans 960 0 0 0 la_data_out[111]
port 302 nsew signal tristate
flabel metal3 s -960 701708 480 701948 0 FreeSans 960 0 0 0 la_data_out[112]
port 303 nsew signal tristate
flabel metal2 s 202206 -960 202318 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 304 nsew signal tristate
flabel metal2 s 570574 703520 570686 704960 0 FreeSans 448 90 0 0 la_data_out[114]
port 305 nsew signal tristate
flabel metal2 s 375442 703520 375554 704960 0 FreeSans 448 90 0 0 la_data_out[115]
port 306 nsew signal tristate
flabel metal2 s 408286 -960 408398 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 307 nsew signal tristate
flabel metal3 s 583520 645268 584960 645508 0 FreeSans 960 0 0 0 la_data_out[117]
port 308 nsew signal tristate
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 la_data_out[118]
port 309 nsew signal tristate
flabel metal3 s 583520 24428 584960 24668 0 FreeSans 960 0 0 0 la_data_out[119]
port 310 nsew signal tristate
flabel metal2 s 452078 703520 452190 704960 0 FreeSans 448 90 0 0 la_data_out[11]
port 311 nsew signal tristate
flabel metal2 s 18666 -960 18778 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 312 nsew signal tristate
flabel metal2 s 184818 703520 184930 704960 0 FreeSans 448 90 0 0 la_data_out[121]
port 313 nsew signal tristate
flabel metal2 s 379306 703520 379418 704960 0 FreeSans 448 90 0 0 la_data_out[122]
port 314 nsew signal tristate
flabel metal3 s -960 229788 480 230028 0 FreeSans 960 0 0 0 la_data_out[123]
port 315 nsew signal tristate
flabel metal3 s 583520 137308 584960 137548 0 FreeSans 960 0 0 0 la_data_out[124]
port 316 nsew signal tristate
flabel metal3 s 583520 480028 584960 480268 0 FreeSans 960 0 0 0 la_data_out[125]
port 317 nsew signal tristate
flabel metal3 s -960 31908 480 32148 0 FreeSans 960 0 0 0 la_data_out[126]
port 318 nsew signal tristate
flabel metal3 s -960 354908 480 355148 0 FreeSans 960 0 0 0 la_data_out[127]
port 319 nsew signal tristate
flabel metal2 s 225390 -960 225502 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 320 nsew signal tristate
flabel metal3 s 583520 40748 584960 40988 0 FreeSans 960 0 0 0 la_data_out[13]
port 321 nsew signal tristate
flabel metal3 s -960 362388 480 362628 0 FreeSans 960 0 0 0 la_data_out[14]
port 322 nsew signal tristate
flabel metal3 s -960 455548 480 455788 0 FreeSans 960 0 0 0 la_data_out[15]
port 323 nsew signal tristate
flabel metal2 s 341310 703520 341422 704960 0 FreeSans 448 90 0 0 la_data_out[16]
port 324 nsew signal tristate
flabel metal3 s 583520 431748 584960 431988 0 FreeSans 960 0 0 0 la_data_out[17]
port 325 nsew signal tristate
flabel metal2 s 110758 -960 110870 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 326 nsew signal tristate
flabel metal2 s 188038 703520 188150 704960 0 FreeSans 448 90 0 0 la_data_out[19]
port 327 nsew signal tristate
flabel metal3 s 583520 93108 584960 93348 0 FreeSans 960 0 0 0 la_data_out[1]
port 328 nsew signal tristate
flabel metal3 s -960 27828 480 28068 0 FreeSans 960 0 0 0 la_data_out[20]
port 329 nsew signal tristate
flabel metal3 s 583520 225708 584960 225948 0 FreeSans 960 0 0 0 la_data_out[21]
port 330 nsew signal tristate
flabel metal3 s 583520 698308 584960 698548 0 FreeSans 960 0 0 0 la_data_out[22]
port 331 nsew signal tristate
flabel metal3 s 583520 229788 584960 230028 0 FreeSans 960 0 0 0 la_data_out[23]
port 332 nsew signal tristate
flabel metal3 s -960 689468 480 689708 0 FreeSans 960 0 0 0 la_data_out[24]
port 333 nsew signal tristate
flabel metal2 s 469466 -960 469578 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 334 nsew signal tristate
flabel metal3 s 583520 467788 584960 468028 0 FreeSans 960 0 0 0 la_data_out[26]
port 335 nsew signal tristate
flabel metal3 s -960 92428 480 92668 0 FreeSans 960 0 0 0 la_data_out[27]
port 336 nsew signal tristate
flabel metal2 s 309110 -960 309222 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 337 nsew signal tristate
flabel metal2 s 305246 -960 305358 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 338 nsew signal tristate
flabel metal2 s 477194 -960 477306 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 339 nsew signal tristate
flabel metal2 s 272402 703520 272514 704960 0 FreeSans 448 90 0 0 la_data_out[30]
port 340 nsew signal tristate
flabel metal3 s -960 237948 480 238188 0 FreeSans 960 0 0 0 la_data_out[31]
port 341 nsew signal tristate
flabel metal3 s -960 217548 480 217788 0 FreeSans 960 0 0 0 la_data_out[32]
port 342 nsew signal tristate
flabel metal3 s 583520 201908 584960 202148 0 FreeSans 960 0 0 0 la_data_out[33]
port 343 nsew signal tristate
flabel metal2 s 316838 -960 316950 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 344 nsew signal tristate
flabel metal3 s -960 322268 480 322508 0 FreeSans 960 0 0 0 la_data_out[35]
port 345 nsew signal tristate
flabel metal2 s 528070 703520 528182 704960 0 FreeSans 448 90 0 0 la_data_out[36]
port 346 nsew signal tristate
flabel metal3 s 583520 8108 584960 8348 0 FreeSans 960 0 0 0 la_data_out[37]
port 347 nsew signal tristate
flabel metal3 s 583520 68628 584960 68868 0 FreeSans 960 0 0 0 la_data_out[38]
port 348 nsew signal tristate
flabel metal3 s 583520 129148 584960 129388 0 FreeSans 960 0 0 0 la_data_out[39]
port 349 nsew signal tristate
flabel metal3 s -960 80188 480 80428 0 FreeSans 960 0 0 0 la_data_out[3]
port 350 nsew signal tristate
flabel metal3 s 583520 346748 584960 346988 0 FreeSans 960 0 0 0 la_data_out[40]
port 351 nsew signal tristate
flabel metal2 s 371578 703520 371690 704960 0 FreeSans 448 90 0 0 la_data_out[41]
port 352 nsew signal tristate
flabel metal2 s 245354 703520 245466 704960 0 FreeSans 448 90 0 0 la_data_out[42]
port 353 nsew signal tristate
flabel metal3 s -960 693548 480 693788 0 FreeSans 960 0 0 0 la_data_out[43]
port 354 nsew signal tristate
flabel metal2 s 465602 -960 465714 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 355 nsew signal tristate
flabel metal2 s 378018 -960 378130 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 356 nsew signal tristate
flabel metal2 s 84998 703520 85110 704960 0 FreeSans 448 90 0 0 la_data_out[46]
port 357 nsew signal tristate
flabel metal3 s -960 628948 480 629188 0 FreeSans 960 0 0 0 la_data_out[47]
port 358 nsew signal tristate
flabel metal2 s 561558 -960 561670 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 359 nsew signal tristate
flabel metal2 s 146178 703520 146290 704960 0 FreeSans 448 90 0 0 la_data_out[49]
port 360 nsew signal tristate
flabel metal2 s 486210 703520 486322 704960 0 FreeSans 448 90 0 0 la_data_out[4]
port 361 nsew signal tristate
flabel metal3 s -960 431068 480 431308 0 FreeSans 960 0 0 0 la_data_out[50]
port 362 nsew signal tristate
flabel metal2 s 370290 -960 370402 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 363 nsew signal tristate
flabel metal3 s -960 84268 480 84508 0 FreeSans 960 0 0 0 la_data_out[52]
port 364 nsew signal tristate
flabel metal2 s 440486 703520 440598 704960 0 FreeSans 448 90 0 0 la_data_out[53]
port 365 nsew signal tristate
flabel metal2 s 397338 -960 397450 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 366 nsew signal tristate
flabel metal3 s -960 201228 480 201468 0 FreeSans 960 0 0 0 la_data_out[55]
port 367 nsew signal tristate
flabel metal2 s 280130 703520 280242 704960 0 FreeSans 448 90 0 0 la_data_out[56]
port 368 nsew signal tristate
flabel metal2 s 47002 703520 47114 704960 0 FreeSans 448 90 0 0 la_data_out[57]
port 369 nsew signal tristate
flabel metal3 s 583520 125068 584960 125308 0 FreeSans 960 0 0 0 la_data_out[58]
port 370 nsew signal tristate
flabel metal3 s 583520 427668 584960 427908 0 FreeSans 960 0 0 0 la_data_out[59]
port 371 nsew signal tristate
flabel metal2 s 354834 -960 354946 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 372 nsew signal tristate
flabel metal3 s -960 645268 480 645508 0 FreeSans 960 0 0 0 la_data_out[60]
port 373 nsew signal tristate
flabel metal3 s -960 411348 480 411588 0 FreeSans 960 0 0 0 la_data_out[61]
port 374 nsew signal tristate
flabel metal2 s 362562 -960 362674 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 375 nsew signal tristate
flabel metal2 s 436622 703520 436734 704960 0 FreeSans 448 90 0 0 la_data_out[63]
port 376 nsew signal tristate
flabel metal3 s -960 273988 480 274228 0 FreeSans 960 0 0 0 la_data_out[64]
port 377 nsew signal tristate
flabel metal2 s 522918 -960 523030 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 378 nsew signal tristate
flabel metal3 s 583520 -52 584960 188 0 FreeSans 960 0 0 0 la_data_out[66]
port 379 nsew signal tristate
flabel metal3 s -960 148868 480 149108 0 FreeSans 960 0 0 0 la_data_out[67]
port 380 nsew signal tristate
flabel metal3 s -960 63868 480 64108 0 FreeSans 960 0 0 0 la_data_out[68]
port 381 nsew signal tristate
flabel metal3 s 583520 181508 584960 181748 0 FreeSans 960 0 0 0 la_data_out[69]
port 382 nsew signal tristate
flabel metal2 s 320702 -960 320814 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 383 nsew signal tristate
flabel metal2 s 473330 -960 473442 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 384 nsew signal tristate
flabel metal3 s -960 48228 480 48468 0 FreeSans 960 0 0 0 la_data_out[71]
port 385 nsew signal tristate
flabel metal2 s 444350 703520 444462 704960 0 FreeSans 448 90 0 0 la_data_out[72]
port 386 nsew signal tristate
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 387 nsew signal tristate
flabel metal2 s 5142 703520 5254 704960 0 FreeSans 448 90 0 0 la_data_out[74]
port 388 nsew signal tristate
flabel metal2 s 400558 -960 400670 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 389 nsew signal tristate
flabel metal3 s -960 669068 480 669308 0 FreeSans 960 0 0 0 la_data_out[76]
port 390 nsew signal tristate
flabel metal3 s 583520 475948 584960 476188 0 FreeSans 960 0 0 0 la_data_out[77]
port 391 nsew signal tristate
flabel metal2 s 332294 -960 332406 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 392 nsew signal tristate
flabel metal3 s 583520 153628 584960 153868 0 FreeSans 960 0 0 0 la_data_out[79]
port 393 nsew signal tristate
flabel metal3 s 583520 44148 584960 44388 0 FreeSans 960 0 0 0 la_data_out[7]
port 394 nsew signal tristate
flabel metal3 s 583520 233868 584960 234108 0 FreeSans 960 0 0 0 la_data_out[80]
port 395 nsew signal tristate
flabel metal3 s -960 572508 480 572748 0 FreeSans 960 0 0 0 la_data_out[81]
port 396 nsew signal tristate
flabel metal2 s 247930 -960 248042 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 397 nsew signal tristate
flabel metal3 s -960 560268 480 560508 0 FreeSans 960 0 0 0 la_data_out[83]
port 398 nsew signal tristate
flabel metal2 s 461738 -960 461850 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 399 nsew signal tristate
flabel metal2 s 517122 703520 517234 704960 0 FreeSans 448 90 0 0 la_data_out[85]
port 400 nsew signal tristate
flabel metal2 s 115910 703520 116022 704960 0 FreeSans 448 90 0 0 la_data_out[86]
port 401 nsew signal tristate
flabel metal2 s 578302 703520 578414 704960 0 FreeSans 448 90 0 0 la_data_out[87]
port 402 nsew signal tristate
flabel metal3 s -960 112828 480 113068 0 FreeSans 960 0 0 0 la_data_out[88]
port 403 nsew signal tristate
flabel metal3 s 583520 76788 584960 77028 0 FreeSans 960 0 0 0 la_data_out[89]
port 404 nsew signal tristate
flabel metal3 s 583520 439908 584960 440148 0 FreeSans 960 0 0 0 la_data_out[8]
port 405 nsew signal tristate
flabel metal2 s 226678 703520 226790 704960 0 FreeSans 448 90 0 0 la_data_out[90]
port 406 nsew signal tristate
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 407 nsew signal tristate
flabel metal2 s 171294 -960 171406 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 408 nsew signal tristate
flabel metal2 s 417302 703520 417414 704960 0 FreeSans 448 90 0 0 la_data_out[93]
port 409 nsew signal tristate
flabel metal2 s 496514 -960 496626 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 410 nsew signal tristate
flabel metal3 s -960 278068 480 278308 0 FreeSans 960 0 0 0 la_data_out[95]
port 411 nsew signal tristate
flabel metal2 s 9006 703520 9118 704960 0 FreeSans 448 90 0 0 la_data_out[96]
port 412 nsew signal tristate
flabel metal2 s 190614 -960 190726 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 413 nsew signal tristate
flabel metal2 s 555118 703520 555230 704960 0 FreeSans 448 90 0 0 la_data_out[98]
port 414 nsew signal tristate
flabel metal2 s 511326 -960 511438 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 415 nsew signal tristate
flabel metal3 s 583520 286228 584960 286468 0 FreeSans 960 0 0 0 la_data_out[9]
port 416 nsew signal tristate
flabel metal2 s 425030 703520 425142 704960 0 FreeSans 448 90 0 0 la_oenb[0]
port 417 nsew signal input
flabel metal3 s -960 209388 480 209628 0 FreeSans 960 0 0 0 la_oenb[100]
port 418 nsew signal input
flabel metal3 s -960 480028 480 480268 0 FreeSans 960 0 0 0 la_oenb[101]
port 419 nsew signal input
flabel metal2 s 297518 -960 297630 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 420 nsew signal input
flabel metal2 s 350970 -960 351082 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 421 nsew signal input
flabel metal2 s 43138 703520 43250 704960 0 FreeSans 448 90 0 0 la_oenb[104]
port 422 nsew signal input
flabel metal3 s 583520 161788 584960 162028 0 FreeSans 960 0 0 0 la_oenb[105]
port 423 nsew signal input
flabel metal2 s 421166 703520 421278 704960 0 FreeSans 448 90 0 0 la_oenb[106]
port 424 nsew signal input
flabel metal2 s 168074 -960 168186 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 425 nsew signal input
flabel metal3 s 583520 471868 584960 472108 0 FreeSans 960 0 0 0 la_oenb[108]
port 426 nsew signal input
flabel metal2 s 177090 703520 177202 704960 0 FreeSans 448 90 0 0 la_oenb[109]
port 427 nsew signal input
flabel metal2 s 513258 703520 513370 704960 0 FreeSans 448 90 0 0 la_oenb[10]
port 428 nsew signal input
flabel metal2 s 142314 703520 142426 704960 0 FreeSans 448 90 0 0 la_oenb[110]
port 429 nsew signal input
flabel metal2 s 35410 703520 35522 704960 0 FreeSans 448 90 0 0 la_oenb[111]
port 430 nsew signal input
flabel metal3 s -960 120308 480 120548 0 FreeSans 960 0 0 0 la_oenb[112]
port 431 nsew signal input
flabel metal2 s 263386 -960 263498 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 432 nsew signal input
flabel metal3 s 583520 596988 584960 597228 0 FreeSans 960 0 0 0 la_oenb[114]
port 433 nsew signal input
flabel metal2 s 481058 -960 481170 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 434 nsew signal input
flabel metal3 s 583520 435828 584960 436068 0 FreeSans 960 0 0 0 la_oenb[116]
port 435 nsew signal input
flabel metal2 s 125570 -960 125682 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 436 nsew signal input
flabel metal2 s 260810 703520 260922 704960 0 FreeSans 448 90 0 0 la_oenb[118]
port 437 nsew signal input
flabel metal3 s -960 44148 480 44388 0 FreeSans 960 0 0 0 la_oenb[119]
port 438 nsew signal input
flabel metal2 s 340022 -960 340134 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 439 nsew signal input
flabel metal2 s 562846 703520 562958 704960 0 FreeSans 448 90 0 0 la_oenb[120]
port 440 nsew signal input
flabel metal3 s -960 378708 480 378948 0 FreeSans 960 0 0 0 la_oenb[121]
port 441 nsew signal input
flabel metal3 s 583520 112828 584960 113068 0 FreeSans 960 0 0 0 la_oenb[122]
port 442 nsew signal input
flabel metal2 s 12870 703520 12982 704960 0 FreeSans 448 90 0 0 la_oenb[123]
port 443 nsew signal input
flabel metal2 s 50866 703520 50978 704960 0 FreeSans 448 90 0 0 la_oenb[124]
port 444 nsew signal input
flabel metal2 s 236338 -960 236450 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 445 nsew signal input
flabel metal2 s 287858 703520 287970 704960 0 FreeSans 448 90 0 0 la_oenb[126]
port 446 nsew signal input
flabel metal3 s 583520 637788 584960 638028 0 FreeSans 960 0 0 0 la_oenb[127]
port 447 nsew signal input
flabel metal3 s 583520 302548 584960 302788 0 FreeSans 960 0 0 0 la_oenb[12]
port 448 nsew signal input
flabel metal3 s -960 318188 480 318428 0 FreeSans 960 0 0 0 la_oenb[13]
port 449 nsew signal input
flabel metal3 s -960 193068 480 193308 0 FreeSans 960 0 0 0 la_oenb[14]
port 450 nsew signal input
flabel metal3 s 583520 246108 584960 246348 0 FreeSans 960 0 0 0 la_oenb[15]
port 451 nsew signal input
flabel metal3 s -960 40068 480 40308 0 FreeSans 960 0 0 0 la_oenb[16]
port 452 nsew signal input
flabel metal2 s 283994 703520 284106 704960 0 FreeSans 448 90 0 0 la_oenb[17]
port 453 nsew signal input
flabel metal3 s -960 152948 480 153188 0 FreeSans 960 0 0 0 la_oenb[18]
port 454 nsew signal input
flabel metal3 s -960 72028 480 72268 0 FreeSans 960 0 0 0 la_oenb[19]
port 455 nsew signal input
flabel metal2 s 186750 -960 186862 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 456 nsew signal input
flabel metal3 s 583520 193748 584960 193988 0 FreeSans 960 0 0 0 la_oenb[20]
port 457 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 458 nsew signal input
flabel metal2 s 194478 -960 194590 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 459 nsew signal input
flabel metal3 s 583520 177428 584960 177668 0 FreeSans 960 0 0 0 la_oenb[23]
port 460 nsew signal input
flabel metal2 s 582166 703520 582278 704960 0 FreeSans 448 90 0 0 la_oenb[24]
port 461 nsew signal input
flabel metal3 s 583520 358988 584960 359228 0 FreeSans 960 0 0 0 la_oenb[25]
port 462 nsew signal input
flabel metal2 s 68254 -960 68366 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 463 nsew signal input
flabel metal3 s 583520 306628 584960 306868 0 FreeSans 960 0 0 0 la_oenb[27]
port 464 nsew signal input
flabel metal3 s -960 15588 480 15828 0 FreeSans 960 0 0 0 la_oenb[28]
port 465 nsew signal input
flabel metal2 s 459806 703520 459918 704960 0 FreeSans 448 90 0 0 la_oenb[29]
port 466 nsew signal input
flabel metal2 s 419878 -960 419990 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 467 nsew signal input
flabel metal3 s 583520 443988 584960 444228 0 FreeSans 960 0 0 0 la_oenb[30]
port 468 nsew signal input
flabel metal2 s 539662 703520 539774 704960 0 FreeSans 448 90 0 0 la_oenb[31]
port 469 nsew signal input
flabel metal3 s -960 23748 480 23988 0 FreeSans 960 0 0 0 la_oenb[32]
port 470 nsew signal input
flabel metal2 s 306534 703520 306646 704960 0 FreeSans 448 90 0 0 la_oenb[33]
port 471 nsew signal input
flabel metal2 s 547390 703520 547502 704960 0 FreeSans 448 90 0 0 la_oenb[34]
port 472 nsew signal input
flabel metal2 s 77270 703520 77382 704960 0 FreeSans 448 90 0 0 la_oenb[35]
port 473 nsew signal input
flabel metal3 s -960 301868 480 302108 0 FreeSans 960 0 0 0 la_oenb[36]
port 474 nsew signal input
flabel metal3 s 583520 116908 584960 117148 0 FreeSans 960 0 0 0 la_oenb[37]
port 475 nsew signal input
flabel metal3 s -960 290308 480 290548 0 FreeSans 960 0 0 0 la_oenb[38]
port 476 nsew signal input
flabel metal3 s 583520 463708 584960 463948 0 FreeSans 960 0 0 0 la_oenb[39]
port 477 nsew signal input
flabel metal2 s 215086 703520 215198 704960 0 FreeSans 448 90 0 0 la_oenb[3]
port 478 nsew signal input
flabel metal2 s 500378 -960 500490 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 479 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 la_oenb[41]
port 480 nsew signal input
flabel metal3 s 583520 532388 584960 532628 0 FreeSans 960 0 0 0 la_oenb[42]
port 481 nsew signal input
flabel metal2 s 490074 703520 490186 704960 0 FreeSans 448 90 0 0 la_oenb[43]
port 482 nsew signal input
flabel metal3 s 583520 681988 584960 682228 0 FreeSans 960 0 0 0 la_oenb[44]
port 483 nsew signal input
flabel metal3 s 583520 16268 584960 16508 0 FreeSans 960 0 0 0 la_oenb[45]
port 484 nsew signal input
flabel metal3 s -960 11508 480 11748 0 FreeSans 960 0 0 0 la_oenb[46]
port 485 nsew signal input
flabel metal2 s 576370 -960 576482 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 486 nsew signal input
flabel metal3 s 583520 108748 584960 108988 0 FreeSans 960 0 0 0 la_oenb[48]
port 487 nsew signal input
flabel metal2 s 117842 -960 117954 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 488 nsew signal input
flabel metal2 s 175158 -960 175270 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 489 nsew signal input
flabel metal3 s 583520 36668 584960 36908 0 FreeSans 960 0 0 0 la_oenb[50]
port 490 nsew signal input
flabel metal3 s 583520 274668 584960 274908 0 FreeSans 960 0 0 0 la_oenb[51]
port 491 nsew signal input
flabel metal3 s 583520 621468 584960 621708 0 FreeSans 960 0 0 0 la_oenb[52]
port 492 nsew signal input
flabel metal2 s 234406 703520 234518 704960 0 FreeSans 448 90 0 0 la_oenb[53]
port 493 nsew signal input
flabel metal2 s 203494 703520 203606 704960 0 FreeSans 448 90 0 0 la_oenb[54]
port 494 nsew signal input
flabel metal2 s 104318 703520 104430 704960 0 FreeSans 448 90 0 0 la_oenb[55]
port 495 nsew signal input
flabel metal2 s 217662 -960 217774 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 496 nsew signal input
flabel metal3 s 583520 690148 584960 690388 0 FreeSans 960 0 0 0 la_oenb[57]
port 497 nsew signal input
flabel metal3 s -960 180828 480 181068 0 FreeSans 960 0 0 0 la_oenb[58]
port 498 nsew signal input
flabel metal2 s 66322 703520 66434 704960 0 FreeSans 448 90 0 0 la_oenb[59]
port 499 nsew signal input
flabel metal3 s -960 52308 480 52548 0 FreeSans 960 0 0 0 la_oenb[5]
port 500 nsew signal input
flabel metal3 s 583520 609228 584960 609468 0 FreeSans 960 0 0 0 la_oenb[60]
port 501 nsew signal input
flabel metal2 s 356122 703520 356234 704960 0 FreeSans 448 90 0 0 la_oenb[61]
port 502 nsew signal input
flabel metal2 s 314262 703520 314374 704960 0 FreeSans 448 90 0 0 la_oenb[62]
port 503 nsew signal input
flabel metal2 s 428894 703520 429006 704960 0 FreeSans 448 90 0 0 la_oenb[63]
port 504 nsew signal input
flabel metal2 s 463670 703520 463782 704960 0 FreeSans 448 90 0 0 la_oenb[64]
port 505 nsew signal input
flabel metal2 s 467534 703520 467646 704960 0 FreeSans 448 90 0 0 la_oenb[65]
port 506 nsew signal input
flabel metal3 s -960 241348 480 241588 0 FreeSans 960 0 0 0 la_oenb[66]
port 507 nsew signal input
flabel metal2 s 249218 703520 249330 704960 0 FreeSans 448 90 0 0 la_oenb[67]
port 508 nsew signal input
flabel metal3 s -960 225708 480 225948 0 FreeSans 960 0 0 0 la_oenb[68]
port 509 nsew signal input
flabel metal2 s 7074 -960 7186 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 510 nsew signal input
flabel metal2 s 572506 -960 572618 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 511 nsew signal input
flabel metal3 s -960 253588 480 253828 0 FreeSans 960 0 0 0 la_oenb[70]
port 512 nsew signal input
flabel metal3 s 583520 197828 584960 198068 0 FreeSans 960 0 0 0 la_oenb[71]
port 513 nsew signal input
flabel metal3 s -960 443308 480 443548 0 FreeSans 960 0 0 0 la_oenb[72]
port 514 nsew signal input
flabel metal3 s 583520 262428 584960 262668 0 FreeSans 960 0 0 0 la_oenb[73]
port 515 nsew signal input
flabel metal3 s -960 584748 480 584988 0 FreeSans 960 0 0 0 la_oenb[74]
port 516 nsew signal input
flabel metal2 s 30258 -960 30370 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 517 nsew signal input
flabel metal3 s -960 261748 480 261988 0 FreeSans 960 0 0 0 la_oenb[76]
port 518 nsew signal input
flabel metal3 s -960 173348 480 173588 0 FreeSans 960 0 0 0 la_oenb[77]
port 519 nsew signal input
flabel metal2 s 242134 703520 242246 704960 0 FreeSans 448 90 0 0 la_oenb[78]
port 520 nsew signal input
flabel metal3 s 583520 4028 584960 4268 0 FreeSans 960 0 0 0 la_oenb[79]
port 521 nsew signal input
flabel metal2 s 278842 -960 278954 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 522 nsew signal input
flabel metal3 s -960 495668 480 495908 0 FreeSans 960 0 0 0 la_oenb[80]
port 523 nsew signal input
flabel metal3 s 583520 528308 584960 528548 0 FreeSans 960 0 0 0 la_oenb[81]
port 524 nsew signal input
flabel metal3 s 583520 669748 584960 669988 0 FreeSans 960 0 0 0 la_oenb[82]
port 525 nsew signal input
flabel metal2 s 565422 -960 565534 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 526 nsew signal input
flabel metal3 s -960 588828 480 589068 0 FreeSans 960 0 0 0 la_oenb[84]
port 527 nsew signal input
flabel metal3 s 583520 141388 584960 141628 0 FreeSans 960 0 0 0 la_oenb[85]
port 528 nsew signal input
flabel metal3 s 583520 633708 584960 633948 0 FreeSans 960 0 0 0 la_oenb[86]
port 529 nsew signal input
flabel metal2 s 153906 703520 154018 704960 0 FreeSans 448 90 0 0 la_oenb[87]
port 530 nsew signal input
flabel metal3 s 583520 540548 584960 540788 0 FreeSans 960 0 0 0 la_oenb[88]
port 531 nsew signal input
flabel metal2 s 549966 -960 550078 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 532 nsew signal input
flabel metal2 s 310398 703520 310510 704960 0 FreeSans 448 90 0 0 la_oenb[8]
port 533 nsew signal input
flabel metal3 s 583520 218228 584960 218468 0 FreeSans 960 0 0 0 la_oenb[90]
port 534 nsew signal input
flabel metal2 s 108182 703520 108294 704960 0 FreeSans 448 90 0 0 la_oenb[91]
port 535 nsew signal input
flabel metal3 s 583520 84948 584960 85188 0 FreeSans 960 0 0 0 la_oenb[92]
port 536 nsew signal input
flabel metal3 s -960 422908 480 423148 0 FreeSans 960 0 0 0 la_oenb[93]
port 537 nsew signal input
flabel metal2 s 91438 -960 91550 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 538 nsew signal input
flabel metal3 s 583520 516748 584960 516988 0 FreeSans 960 0 0 0 la_oenb[95]
port 539 nsew signal input
flabel metal2 s 404422 -960 404534 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 540 nsew signal input
flabel metal3 s -960 221628 480 221868 0 FreeSans 960 0 0 0 la_oenb[97]
port 541 nsew signal input
flabel metal2 s 182886 -960 182998 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 542 nsew signal input
flabel metal3 s -960 294388 480 294628 0 FreeSans 960 0 0 0 la_oenb[99]
port 543 nsew signal input
flabel metal3 s -960 616708 480 616948 0 FreeSans 960 0 0 0 la_oenb[9]
port 544 nsew signal input
flabel metal2 s 318126 703520 318238 704960 0 FreeSans 448 90 0 0 user_clock2
port 545 nsew signal input
flabel metal3 s 583520 702388 584960 702628 0 FreeSans 960 0 0 0 user_irq[0]
port 546 nsew signal tristate
flabel metal3 s -960 596988 480 597228 0 FreeSans 960 0 0 0 user_irq[1]
port 547 nsew signal tristate
flabel metal3 s -960 660908 480 661148 0 FreeSans 960 0 0 0 user_irq[2]
port 548 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 549 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 550 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 551 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 552 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 553 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 554 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 555 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 556 nsew ground bidirectional
flabel metal3 s 583520 258348 584960 258588 0 FreeSans 960 0 0 0 wb_clk_i
port 557 nsew signal input
flabel metal3 s -960 350828 480 351068 0 FreeSans 960 0 0 0 wb_rst_i
port 558 nsew signal input
flabel metal3 s 583520 383468 584960 383708 0 FreeSans 960 0 0 0 wbs_ack_o
port 559 nsew signal tristate
flabel metal2 s 199630 703520 199742 704960 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 560 nsew signal input
flabel metal2 s 54730 703520 54842 704960 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 561 nsew signal input
flabel metal3 s -960 471868 480 472108 0 FreeSans 960 0 0 0 wbs_adr_i[11]
port 562 nsew signal input
flabel metal2 s 64390 -960 64502 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 563 nsew signal input
flabel metal2 s 389610 -960 389722 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 564 nsew signal input
flabel metal3 s 583520 657508 584960 657748 0 FreeSans 960 0 0 0 wbs_adr_i[14]
port 565 nsew signal input
flabel metal3 s 583520 613308 584960 613548 0 FreeSans 960 0 0 0 wbs_adr_i[15]
port 566 nsew signal input
flabel metal2 s 443062 -960 443174 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 567 nsew signal input
flabel metal3 s 583520 556868 584960 557108 0 FreeSans 960 0 0 0 wbs_adr_i[17]
port 568 nsew signal input
flabel metal3 s 583520 343348 584960 343588 0 FreeSans 960 0 0 0 wbs_adr_i[18]
port 569 nsew signal input
flabel metal3 s 583520 89028 584960 89268 0 FreeSans 960 0 0 0 wbs_adr_i[19]
port 570 nsew signal input
flabel metal2 s 207358 703520 207470 704960 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 571 nsew signal input
flabel metal2 s 406354 703520 406466 704960 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 572 nsew signal input
flabel metal2 s 393474 -960 393586 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 573 nsew signal input
flabel metal2 s 557694 -960 557806 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 574 nsew signal input
flabel metal3 s 583520 278748 584960 278988 0 FreeSans 960 0 0 0 wbs_adr_i[23]
port 575 nsew signal input
flabel metal3 s -960 556188 480 556428 0 FreeSans 960 0 0 0 wbs_adr_i[24]
port 576 nsew signal input
flabel metal2 s 374154 -960 374266 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 577 nsew signal input
flabel metal2 s 72118 -960 72230 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 578 nsew signal input
flabel metal3 s -960 19668 480 19908 0 FreeSans 960 0 0 0 wbs_adr_i[27]
port 579 nsew signal input
flabel metal3 s 583520 524228 584960 524468 0 FreeSans 960 0 0 0 wbs_adr_i[28]
port 580 nsew signal input
flabel metal2 s 497802 703520 497914 704960 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 581 nsew signal input
flabel metal2 s 267250 -960 267362 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 582 nsew signal input
flabel metal2 s 333582 703520 333694 704960 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 583 nsew signal input
flabel metal3 s 583520 403868 584960 404108 0 FreeSans 960 0 0 0 wbs_adr_i[31]
port 584 nsew signal input
flabel metal2 s 530646 -960 530758 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 585 nsew signal input
flabel metal2 s 321990 703520 322102 704960 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 586 nsew signal input
flabel metal3 s -960 108748 480 108988 0 FreeSans 960 0 0 0 wbs_adr_i[5]
port 587 nsew signal input
flabel metal2 s 213798 -960 213910 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 588 nsew signal input
flabel metal2 s 34122 -960 34234 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 589 nsew signal input
flabel metal3 s 583520 97188 584960 97428 0 FreeSans 960 0 0 0 wbs_adr_i[8]
port 590 nsew signal input
flabel metal3 s 583520 290308 584960 290548 0 FreeSans 960 0 0 0 wbs_adr_i[9]
port 591 nsew signal input
flabel metal2 s 31546 703520 31658 704960 0 FreeSans 448 90 0 0 wbs_cyc_i
port 592 nsew signal input
flabel metal2 s 574438 703520 574550 704960 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 593 nsew signal input
flabel metal3 s -960 358988 480 359228 0 FreeSans 960 0 0 0 wbs_dat_i[10]
port 594 nsew signal input
flabel metal3 s -960 407268 480 407508 0 FreeSans 960 0 0 0 wbs_dat_i[11]
port 595 nsew signal input
flabel metal3 s -960 390948 480 391188 0 FreeSans 960 0 0 0 wbs_dat_i[12]
port 596 nsew signal input
flabel metal2 s 26394 -960 26506 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 597 nsew signal input
flabel metal2 s 144890 -960 145002 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 598 nsew signal input
flabel metal3 s 583520 456228 584960 456468 0 FreeSans 960 0 0 0 wbs_dat_i[15]
port 599 nsew signal input
flabel metal2 s 385746 -960 385858 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 600 nsew signal input
flabel metal2 s 291722 703520 291834 704960 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 601 nsew signal input
flabel metal2 s 455942 703520 456054 704960 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 602 nsew signal input
flabel metal3 s -960 576588 480 576828 0 FreeSans 960 0 0 0 wbs_dat_i[19]
port 603 nsew signal input
flabel metal2 s 103030 -960 103142 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 604 nsew signal input
flabel metal3 s 583520 508588 584960 508828 0 FreeSans 960 0 0 0 wbs_dat_i[20]
port 605 nsew signal input
flabel metal2 s 482346 703520 482458 704960 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 606 nsew signal input
flabel metal3 s -960 265828 480 266068 0 FreeSans 960 0 0 0 wbs_dat_i[22]
port 607 nsew signal input
flabel metal3 s 583520 629628 584960 629868 0 FreeSans 960 0 0 0 wbs_dat_i[23]
port 608 nsew signal input
flabel metal3 s 583520 310708 584960 310948 0 FreeSans 960 0 0 0 wbs_dat_i[24]
port 609 nsew signal input
flabel metal2 s 457874 -960 457986 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 610 nsew signal input
flabel metal2 s 410218 703520 410330 704960 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 611 nsew signal input
flabel metal2 s 19954 703520 20066 704960 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 612 nsew signal input
flabel metal2 s 206070 -960 206182 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 613 nsew signal input
flabel metal3 s 583520 496348 584960 496588 0 FreeSans 960 0 0 0 wbs_dat_i[29]
port 614 nsew signal input
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 615 nsew signal input
flabel metal3 s 583520 282828 584960 283068 0 FreeSans 960 0 0 0 wbs_dat_i[30]
port 616 nsew signal input
flabel metal3 s -960 249508 480 249748 0 FreeSans 960 0 0 0 wbs_dat_i[31]
port 617 nsew signal input
flabel metal3 s 583520 101268 584960 101508 0 FreeSans 960 0 0 0 wbs_dat_i[3]
port 618 nsew signal input
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 619 nsew signal input
flabel metal2 s 324566 -960 324678 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 620 nsew signal input
flabel metal3 s -960 3348 480 3588 0 FreeSans 960 0 0 0 wbs_dat_i[6]
port 621 nsew signal input
flabel metal2 s 398626 703520 398738 704960 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 622 nsew signal input
flabel metal3 s 583520 686068 584960 686308 0 FreeSans 960 0 0 0 wbs_dat_i[8]
port 623 nsew signal input
flabel metal3 s 583520 104668 584960 104908 0 FreeSans 960 0 0 0 wbs_dat_i[9]
port 624 nsew signal input
flabel metal2 s 53442 -960 53554 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 625 nsew signal tristate
flabel metal3 s 583520 460308 584960 460548 0 FreeSans 960 0 0 0 wbs_dat_o[10]
port 626 nsew signal tristate
flabel metal2 s 14802 -960 14914 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 627 nsew signal tristate
flabel metal3 s 583520 694228 584960 694468 0 FreeSans 960 0 0 0 wbs_dat_o[12]
port 628 nsew signal tristate
flabel metal2 s 383170 703520 383282 704960 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 629 nsew signal tristate
flabel metal3 s 583520 145468 584960 145708 0 FreeSans 960 0 0 0 wbs_dat_o[14]
port 630 nsew signal tristate
flabel metal2 s 363850 703520 363962 704960 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 631 nsew signal tristate
flabel metal3 s -960 116908 480 117148 0 FreeSans 960 0 0 0 wbs_dat_o[16]
port 632 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 wbs_dat_o[17]
port 633 nsew signal tristate
flabel metal2 s 435334 -960 435446 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 634 nsew signal tristate
flabel metal2 s -10 -960 102 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 635 nsew signal tristate
flabel metal2 s 508106 -960 508218 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 636 nsew signal tristate
flabel metal3 s -960 257668 480 257908 0 FreeSans 960 0 0 0 wbs_dat_o[20]
port 637 nsew signal tristate
flabel metal3 s -960 524228 480 524468 0 FreeSans 960 0 0 0 wbs_dat_o[21]
port 638 nsew signal tristate
flabel metal2 s 92726 703520 92838 704960 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 639 nsew signal tristate
flabel metal3 s -960 169268 480 169508 0 FreeSans 960 0 0 0 wbs_dat_o[23]
port 640 nsew signal tristate
flabel metal2 s 133298 -960 133410 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 641 nsew signal tristate
flabel metal2 s 49578 -960 49690 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 642 nsew signal tristate
flabel metal2 s 256946 703520 257058 704960 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 643 nsew signal tristate
flabel metal2 s 112046 703520 112158 704960 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 644 nsew signal tristate
flabel metal2 s 347106 -960 347218 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 645 nsew signal tristate
flabel metal2 s 367714 703520 367826 704960 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 646 nsew signal tristate
flabel metal3 s 583520 242028 584960 242268 0 FreeSans 960 0 0 0 wbs_dat_o[2]
port 647 nsew signal tristate
flabel metal3 s -960 403188 480 403428 0 FreeSans 960 0 0 0 wbs_dat_o[30]
port 648 nsew signal tristate
flabel metal3 s 583520 569108 584960 569348 0 FreeSans 960 0 0 0 wbs_dat_o[31]
port 649 nsew signal tristate
flabel metal2 s 141026 -960 141138 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 650 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 651 nsew signal tristate
flabel metal3 s -960 35988 480 36228 0 FreeSans 960 0 0 0 wbs_dat_o[5]
port 652 nsew signal tristate
flabel metal3 s 583520 544628 584960 544868 0 FreeSans 960 0 0 0 wbs_dat_o[6]
port 653 nsew signal tristate
flabel metal2 s 381882 -960 381994 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 654 nsew signal tristate
flabel metal2 s 359986 703520 360098 704960 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 655 nsew signal tristate
flabel metal2 s 352902 703520 353014 704960 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 656 nsew signal tristate
flabel metal3 s -960 600388 480 600628 0 FreeSans 960 0 0 0 wbs_sel_i[0]
port 657 nsew signal input
flabel metal2 s 16090 703520 16202 704960 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 658 nsew signal input
flabel metal2 s 454654 -960 454766 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 659 nsew signal input
flabel metal3 s -960 140708 480 140948 0 FreeSans 960 0 0 0 wbs_sel_i[3]
port 660 nsew signal input
flabel metal3 s -960 543948 480 544188 0 FreeSans 960 0 0 0 wbs_stb_i
port 661 nsew signal input
flabel metal3 s 583520 371228 584960 371468 0 FreeSans 960 0 0 0 wbs_we_i
port 662 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
